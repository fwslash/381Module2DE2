// nios2_system.v

// Generated using ACDS version 13.0sp1 232 at 2014.11.12.17:22:29

`timescale 1 ps / 1 ps
module nios2_system (
		input  wire        clk_clk,                                         //                                       clk.clk
		input  wire        reset_reset_n,                                   //                                     reset.reset_n
		output wire [11:0] sdram_wire_addr,                                 //                                sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                                   //                                          .ba
		output wire        sdram_wire_cas_n,                                //                                          .cas_n
		output wire        sdram_wire_cke,                                  //                                          .cke
		output wire        sdram_wire_cs_n,                                 //                                          .cs_n
		inout  wire [15:0] sdram_wire_dq,                                   //                                          .dq
		output wire [1:0]  sdram_wire_dqm,                                  //                                          .dqm
		output wire        sdram_wire_ras_n,                                //                                          .ras_n
		output wire        sdram_wire_we_n,                                 //                                          .we_n
		output wire [7:0]  ledg_export,                                     //                                      ledg.export
		output wire [17:0] ledr_export,                                     //                                      ledr.export
		input  wire [17:0] switches_export,                                 //                                  switches.export
		input  wire [3:0]  keys_export,                                     //                                      keys.export
		inout  wire [7:0]  lcd_data_DATA,                                   //                                  lcd_data.DATA
		output wire        lcd_data_ON,                                     //                                          .ON
		output wire        lcd_data_BLON,                                   //                                          .BLON
		output wire        lcd_data_EN,                                     //                                          .EN
		output wire        lcd_data_RS,                                     //                                          .RS
		output wire        lcd_data_RW,                                     //                                          .RW
		output wire        video_vga_controller_0_external_interface_CLK,   // video_vga_controller_0_external_interface.CLK
		output wire        video_vga_controller_0_external_interface_HS,    //                                          .HS
		output wire        video_vga_controller_0_external_interface_VS,    //                                          .VS
		output wire        video_vga_controller_0_external_interface_BLANK, //                                          .BLANK
		output wire        video_vga_controller_0_external_interface_SYNC,  //                                          .SYNC
		output wire [9:0]  video_vga_controller_0_external_interface_R,     //                                          .R
		output wire [9:0]  video_vga_controller_0_external_interface_G,     //                                          .G
		output wire [9:0]  video_vga_controller_0_external_interface_B,     //                                          .B
		inout  wire        sdcard_b_SD_cmd,                                 //                                    sdcard.b_SD_cmd
		inout  wire        sdcard_b_SD_dat,                                 //                                          .b_SD_dat
		inout  wire        sdcard_b_SD_dat3,                                //                                          .b_SD_dat3
		output wire        sdcard_o_SD_clock,                               //                                          .o_SD_clock
		inout  wire        ps2_peri_CLK,                                    //                                  ps2_peri.CLK
		inout  wire        ps2_peri_DAT,                                    //                                          .DAT
		inout  wire [15:0] sram_0_external_interface_DQ,                    //                 sram_0_external_interface.DQ
		output wire [17:0] sram_0_external_interface_ADDR,                  //                                          .ADDR
		output wire        sram_0_external_interface_LB_N,                  //                                          .LB_N
		output wire        sram_0_external_interface_UB_N,                  //                                          .UB_N
		output wire        sram_0_external_interface_CE_N,                  //                                          .CE_N
		output wire        sram_0_external_interface_OE_N,                  //                                          .OE_N
		output wire        sram_0_external_interface_WE_N,                  //                                          .WE_N
		input  wire        audio_ADCDAT,                                    //                                     audio.ADCDAT
		input  wire        audio_ADCLRCK,                                   //                                          .ADCLRCK
		input  wire        audio_BCLK,                                      //                                          .BCLK
		output wire        audio_DACDAT,                                    //                                          .DACDAT
		input  wire        audio_DACLRCK,                                   //                                          .DACLRCK
		output wire        sdram_clk_clk,                                   //                                 sdram_clk.clk
		input  wire        audio_secondary_clk,                             //                           audio_secondary.clk
		output wire        audio_clk_clk,                                   //                                 audio_clk.clk
		inout  wire        av_config_SDAT,                                  //                                 av_config.SDAT
		output wire        av_config_SCLK,                                  //                                          .SCLK
		input  wire        usb_INT1,                                        //                                       usb.INT1
		inout  wire [15:0] usb_DATA,                                        //                                          .DATA
		output wire        usb_RST_N,                                       //                                          .RST_N
		output wire [1:0]  usb_ADDR,                                        //                                          .ADDR
		output wire        usb_CS_N,                                        //                                          .CS_N
		output wire        usb_RD_N,                                        //                                          .RD_N
		output wire        usb_WR_N,                                        //                                          .WR_N
		input  wire        usb_INT0                                         //                                          .INT0
	);

	wire          clocks_sys_clk_clk;                                                                                                               // clocks:sys_clk -> [Altera_UP_SD_Card_Avalon_Interface_0:i_clock, Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:clk, Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:clk, Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, JTAG:clk, JTAG_avalon_jtag_slave_translator:clk, JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, LEDG:clk, LEDG_s1_translator:clk, LEDG_s1_translator_avalon_universal_slave_0_agent:clk, LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, LEDR:clk, LEDR_s1_translator:clk, LEDR_s1_translator_avalon_universal_slave_0_agent:clk, LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, addr_router:clk, addr_router_001:clk, addr_router_002:clk, audio_0:clk, audio_0_avalon_audio_slave_translator:clk, audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:clk, audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, audio_and_video_config_0:clk, audio_and_video_config_0_avalon_av_config_slave_translator:clk, audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:clk, audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, burst_adapter:clk, burst_adapter_001:clk, burst_adapter_002:clk, burst_adapter_003:clk, character_lcd_0:clk, character_lcd_0_avalon_lcd_slave_translator:clk, character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:clk, character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_demux_002:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, cmd_xbar_mux_002:clk, cmd_xbar_mux_003:clk, cmd_xbar_mux_004:clk, cmd_xbar_mux_005:clk, cmd_xbar_mux_006:clk, cmd_xbar_mux_007:clk, cmd_xbar_mux_008:clk, cmd_xbar_mux_009:clk, cmd_xbar_mux_010:clk, cmd_xbar_mux_016:clk, cmd_xbar_mux_018:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, id_router_006:clk, id_router_007:clk, id_router_008:clk, id_router_009:clk, id_router_010:clk, id_router_011:clk, id_router_012:clk, id_router_013:clk, id_router_014:clk, id_router_015:clk, id_router_016:clk, id_router_017:clk, id_router_018:clk, irq_mapper:clk, key:clk, key_s1_translator:clk, key_s1_translator_avalon_universal_slave_0_agent:clk, key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, limiter:clk, limiter_001:clk, limiter_002:clk, nios2_system:clk, nios2_system_data_master_translator:clk, nios2_system_data_master_translator_avalon_universal_master_0_agent:clk, nios2_system_instruction_master_translator:clk, nios2_system_instruction_master_translator_avalon_universal_master_0_agent:clk, nios2_system_jtag_debug_module_translator:clk, nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, onchip:clk, onchip_s1_translator:clk, onchip_s1_translator_avalon_universal_slave_0_agent:clk, onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, ps2_0:clk, ps2_0_avalon_ps2_slave_translator:clk, ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:clk, ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_demux_009:clk, rsp_xbar_demux_010:clk, rsp_xbar_demux_011:clk, rsp_xbar_demux_012:clk, rsp_xbar_demux_013:clk, rsp_xbar_demux_014:clk, rsp_xbar_demux_015:clk, rsp_xbar_demux_016:clk, rsp_xbar_demux_017:clk, rsp_xbar_demux_018:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rsp_xbar_mux_002:clk, rst_controller:clk, sdcard_timer:clk, sdcard_timer_s1_translator:clk, sdcard_timer_s1_translator_avalon_universal_slave_0_agent:clk, sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sdram:clk, sdram_s1_translator:clk, sdram_s1_translator_avalon_universal_slave_0_agent:clk, sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sram_0:clk, sram_0_avalon_sram_slave_translator:clk, sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:clk, sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, switches:clk, switches_s1_translator:clk, switches_s1_translator_avalon_universal_slave_0_agent:clk, switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, usb_0:clk, usb_0_avalon_usb_slave_translator:clk, usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:clk, usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, video_alpha_blender_0:clk, video_character_buffer_with_dma_0:clk, video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator:clk, video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:clk, video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, video_character_buffer_with_dma_0_avalon_char_control_slave_translator:clk, video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:clk, video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, video_dual_clock_buffer_0:clk_stream_in, video_pixel_buffer_dma:clk, video_pixel_buffer_dma_avalon_control_slave_translator:clk, video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:clk, video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, video_pixel_buffer_dma_avalon_pixel_dma_master_translator:clk, video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:clk, video_rgb_resampler_0:clk, video_scaler_0:clk, width_adapter:clk, width_adapter_001:clk, width_adapter_002:clk, width_adapter_003:clk, width_adapter_004:clk, width_adapter_005:clk, width_adapter_006:clk, width_adapter_007:clk, width_adapter_008:clk, width_adapter_009:clk, width_adapter_010:clk, width_adapter_011:clk]
	wire          video_pixel_buffer_dma_avalon_pixel_source_endofpacket;                                                                           // video_pixel_buffer_dma:stream_endofpacket -> video_rgb_resampler_0:stream_in_endofpacket
	wire          video_pixel_buffer_dma_avalon_pixel_source_valid;                                                                                 // video_pixel_buffer_dma:stream_valid -> video_rgb_resampler_0:stream_in_valid
	wire          video_pixel_buffer_dma_avalon_pixel_source_startofpacket;                                                                         // video_pixel_buffer_dma:stream_startofpacket -> video_rgb_resampler_0:stream_in_startofpacket
	wire   [15:0] video_pixel_buffer_dma_avalon_pixel_source_data;                                                                                  // video_pixel_buffer_dma:stream_data -> video_rgb_resampler_0:stream_in_data
	wire          video_pixel_buffer_dma_avalon_pixel_source_ready;                                                                                 // video_rgb_resampler_0:stream_in_ready -> video_pixel_buffer_dma:stream_ready
	wire          clocks_vga_clk_clk;                                                                                                               // clocks:VGA_CLK -> [rst_controller_002:clk, video_dual_clock_buffer_0:clk_stream_out, video_vga_controller_0:clk]
	wire          video_character_buffer_with_dma_0_avalon_char_source_endofpacket;                                                                 // video_character_buffer_with_dma_0:stream_endofpacket -> video_alpha_blender_0:foreground_endofpacket
	wire          video_character_buffer_with_dma_0_avalon_char_source_valid;                                                                       // video_character_buffer_with_dma_0:stream_valid -> video_alpha_blender_0:foreground_valid
	wire          video_character_buffer_with_dma_0_avalon_char_source_startofpacket;                                                               // video_character_buffer_with_dma_0:stream_startofpacket -> video_alpha_blender_0:foreground_startofpacket
	wire   [39:0] video_character_buffer_with_dma_0_avalon_char_source_data;                                                                        // video_character_buffer_with_dma_0:stream_data -> video_alpha_blender_0:foreground_data
	wire          video_character_buffer_with_dma_0_avalon_char_source_ready;                                                                       // video_alpha_blender_0:foreground_ready -> video_character_buffer_with_dma_0:stream_ready
	wire          video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket;                                                                    // video_dual_clock_buffer_0:stream_out_endofpacket -> video_vga_controller_0:endofpacket
	wire          video_dual_clock_buffer_0_avalon_dc_buffer_source_valid;                                                                          // video_dual_clock_buffer_0:stream_out_valid -> video_vga_controller_0:valid
	wire          video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket;                                                                  // video_dual_clock_buffer_0:stream_out_startofpacket -> video_vga_controller_0:startofpacket
	wire   [29:0] video_dual_clock_buffer_0_avalon_dc_buffer_source_data;                                                                           // video_dual_clock_buffer_0:stream_out_data -> video_vga_controller_0:data
	wire          video_dual_clock_buffer_0_avalon_dc_buffer_source_ready;                                                                          // video_vga_controller_0:ready -> video_dual_clock_buffer_0:stream_out_ready
	wire          video_scaler_0_avalon_scaler_source_endofpacket;                                                                                  // video_scaler_0:stream_out_endofpacket -> video_alpha_blender_0:background_endofpacket
	wire          video_scaler_0_avalon_scaler_source_valid;                                                                                        // video_scaler_0:stream_out_valid -> video_alpha_blender_0:background_valid
	wire          video_scaler_0_avalon_scaler_source_startofpacket;                                                                                // video_scaler_0:stream_out_startofpacket -> video_alpha_blender_0:background_startofpacket
	wire   [29:0] video_scaler_0_avalon_scaler_source_data;                                                                                         // video_scaler_0:stream_out_data -> video_alpha_blender_0:background_data
	wire          video_scaler_0_avalon_scaler_source_ready;                                                                                        // video_alpha_blender_0:background_ready -> video_scaler_0:stream_out_ready
	wire          video_rgb_resampler_0_avalon_rgb_source_endofpacket;                                                                              // video_rgb_resampler_0:stream_out_endofpacket -> video_scaler_0:stream_in_endofpacket
	wire          video_rgb_resampler_0_avalon_rgb_source_valid;                                                                                    // video_rgb_resampler_0:stream_out_valid -> video_scaler_0:stream_in_valid
	wire          video_rgb_resampler_0_avalon_rgb_source_startofpacket;                                                                            // video_rgb_resampler_0:stream_out_startofpacket -> video_scaler_0:stream_in_startofpacket
	wire   [29:0] video_rgb_resampler_0_avalon_rgb_source_data;                                                                                     // video_rgb_resampler_0:stream_out_data -> video_scaler_0:stream_in_data
	wire          video_rgb_resampler_0_avalon_rgb_source_ready;                                                                                    // video_scaler_0:stream_in_ready -> video_rgb_resampler_0:stream_out_ready
	wire          video_alpha_blender_0_avalon_blended_source_endofpacket;                                                                          // video_alpha_blender_0:output_endofpacket -> video_dual_clock_buffer_0:stream_in_endofpacket
	wire          video_alpha_blender_0_avalon_blended_source_valid;                                                                                // video_alpha_blender_0:output_valid -> video_dual_clock_buffer_0:stream_in_valid
	wire          video_alpha_blender_0_avalon_blended_source_startofpacket;                                                                        // video_alpha_blender_0:output_startofpacket -> video_dual_clock_buffer_0:stream_in_startofpacket
	wire   [29:0] video_alpha_blender_0_avalon_blended_source_data;                                                                                 // video_alpha_blender_0:output_data -> video_dual_clock_buffer_0:stream_in_data
	wire          video_alpha_blender_0_avalon_blended_source_ready;                                                                                // video_dual_clock_buffer_0:stream_in_ready -> video_alpha_blender_0:output_ready
	wire          nios2_system_instruction_master_waitrequest;                                                                                      // nios2_system_instruction_master_translator:av_waitrequest -> nios2_system:i_waitrequest
	wire   [24:0] nios2_system_instruction_master_address;                                                                                          // nios2_system:i_address -> nios2_system_instruction_master_translator:av_address
	wire          nios2_system_instruction_master_read;                                                                                             // nios2_system:i_read -> nios2_system_instruction_master_translator:av_read
	wire   [31:0] nios2_system_instruction_master_readdata;                                                                                         // nios2_system_instruction_master_translator:av_readdata -> nios2_system:i_readdata
	wire          nios2_system_instruction_master_readdatavalid;                                                                                    // nios2_system_instruction_master_translator:av_readdatavalid -> nios2_system:i_readdatavalid
	wire          nios2_system_data_master_waitrequest;                                                                                             // nios2_system_data_master_translator:av_waitrequest -> nios2_system:d_waitrequest
	wire   [31:0] nios2_system_data_master_writedata;                                                                                               // nios2_system:d_writedata -> nios2_system_data_master_translator:av_writedata
	wire   [24:0] nios2_system_data_master_address;                                                                                                 // nios2_system:d_address -> nios2_system_data_master_translator:av_address
	wire          nios2_system_data_master_write;                                                                                                   // nios2_system:d_write -> nios2_system_data_master_translator:av_write
	wire          nios2_system_data_master_read;                                                                                                    // nios2_system:d_read -> nios2_system_data_master_translator:av_read
	wire   [31:0] nios2_system_data_master_readdata;                                                                                                // nios2_system_data_master_translator:av_readdata -> nios2_system:d_readdata
	wire          nios2_system_data_master_debugaccess;                                                                                             // nios2_system:jtag_debug_module_debugaccess_to_roms -> nios2_system_data_master_translator:av_debugaccess
	wire          nios2_system_data_master_readdatavalid;                                                                                           // nios2_system_data_master_translator:av_readdatavalid -> nios2_system:d_readdatavalid
	wire    [3:0] nios2_system_data_master_byteenable;                                                                                              // nios2_system:d_byteenable -> nios2_system_data_master_translator:av_byteenable
	wire          video_pixel_buffer_dma_avalon_pixel_dma_master_waitrequest;                                                                       // video_pixel_buffer_dma_avalon_pixel_dma_master_translator:av_waitrequest -> video_pixel_buffer_dma:master_waitrequest
	wire   [31:0] video_pixel_buffer_dma_avalon_pixel_dma_master_address;                                                                           // video_pixel_buffer_dma:master_address -> video_pixel_buffer_dma_avalon_pixel_dma_master_translator:av_address
	wire          video_pixel_buffer_dma_avalon_pixel_dma_master_lock;                                                                              // video_pixel_buffer_dma:master_arbiterlock -> video_pixel_buffer_dma_avalon_pixel_dma_master_translator:av_lock
	wire          video_pixel_buffer_dma_avalon_pixel_dma_master_read;                                                                              // video_pixel_buffer_dma:master_read -> video_pixel_buffer_dma_avalon_pixel_dma_master_translator:av_read
	wire   [15:0] video_pixel_buffer_dma_avalon_pixel_dma_master_readdata;                                                                          // video_pixel_buffer_dma_avalon_pixel_dma_master_translator:av_readdata -> video_pixel_buffer_dma:master_readdata
	wire          video_pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid;                                                                     // video_pixel_buffer_dma_avalon_pixel_dma_master_translator:av_readdatavalid -> video_pixel_buffer_dma:master_readdatavalid
	wire          nios2_system_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                                                        // nios2_system:jtag_debug_module_waitrequest -> nios2_system_jtag_debug_module_translator:av_waitrequest
	wire   [31:0] nios2_system_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                                          // nios2_system_jtag_debug_module_translator:av_writedata -> nios2_system:jtag_debug_module_writedata
	wire    [8:0] nios2_system_jtag_debug_module_translator_avalon_anti_slave_0_address;                                                            // nios2_system_jtag_debug_module_translator:av_address -> nios2_system:jtag_debug_module_address
	wire          nios2_system_jtag_debug_module_translator_avalon_anti_slave_0_write;                                                              // nios2_system_jtag_debug_module_translator:av_write -> nios2_system:jtag_debug_module_write
	wire          nios2_system_jtag_debug_module_translator_avalon_anti_slave_0_read;                                                               // nios2_system_jtag_debug_module_translator:av_read -> nios2_system:jtag_debug_module_read
	wire   [31:0] nios2_system_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                                           // nios2_system:jtag_debug_module_readdata -> nios2_system_jtag_debug_module_translator:av_readdata
	wire          nios2_system_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                                        // nios2_system_jtag_debug_module_translator:av_debugaccess -> nios2_system:jtag_debug_module_debugaccess
	wire    [3:0] nios2_system_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                                         // nios2_system_jtag_debug_module_translator:av_byteenable -> nios2_system:jtag_debug_module_byteenable
	wire   [31:0] onchip_s1_translator_avalon_anti_slave_0_writedata;                                                                               // onchip_s1_translator:av_writedata -> onchip:writedata
	wire    [9:0] onchip_s1_translator_avalon_anti_slave_0_address;                                                                                 // onchip_s1_translator:av_address -> onchip:address
	wire          onchip_s1_translator_avalon_anti_slave_0_chipselect;                                                                              // onchip_s1_translator:av_chipselect -> onchip:chipselect
	wire          onchip_s1_translator_avalon_anti_slave_0_clken;                                                                                   // onchip_s1_translator:av_clken -> onchip:clken
	wire          onchip_s1_translator_avalon_anti_slave_0_write;                                                                                   // onchip_s1_translator:av_write -> onchip:write
	wire   [31:0] onchip_s1_translator_avalon_anti_slave_0_readdata;                                                                                // onchip:readdata -> onchip_s1_translator:av_readdata
	wire    [3:0] onchip_s1_translator_avalon_anti_slave_0_byteenable;                                                                              // onchip_s1_translator:av_byteenable -> onchip:byteenable
	wire          sdram_s1_translator_avalon_anti_slave_0_waitrequest;                                                                              // sdram:za_waitrequest -> sdram_s1_translator:av_waitrequest
	wire   [15:0] sdram_s1_translator_avalon_anti_slave_0_writedata;                                                                                // sdram_s1_translator:av_writedata -> sdram:az_data
	wire   [21:0] sdram_s1_translator_avalon_anti_slave_0_address;                                                                                  // sdram_s1_translator:av_address -> sdram:az_addr
	wire          sdram_s1_translator_avalon_anti_slave_0_chipselect;                                                                               // sdram_s1_translator:av_chipselect -> sdram:az_cs
	wire          sdram_s1_translator_avalon_anti_slave_0_write;                                                                                    // sdram_s1_translator:av_write -> sdram:az_wr_n
	wire          sdram_s1_translator_avalon_anti_slave_0_read;                                                                                     // sdram_s1_translator:av_read -> sdram:az_rd_n
	wire   [15:0] sdram_s1_translator_avalon_anti_slave_0_readdata;                                                                                 // sdram:za_data -> sdram_s1_translator:av_readdata
	wire          sdram_s1_translator_avalon_anti_slave_0_readdatavalid;                                                                            // sdram:za_valid -> sdram_s1_translator:av_readdatavalid
	wire    [1:0] sdram_s1_translator_avalon_anti_slave_0_byteenable;                                                                               // sdram_s1_translator:av_byteenable -> sdram:az_be_n
	wire   [31:0] ledg_s1_translator_avalon_anti_slave_0_writedata;                                                                                 // LEDG_s1_translator:av_writedata -> LEDG:writedata
	wire    [1:0] ledg_s1_translator_avalon_anti_slave_0_address;                                                                                   // LEDG_s1_translator:av_address -> LEDG:address
	wire          ledg_s1_translator_avalon_anti_slave_0_chipselect;                                                                                // LEDG_s1_translator:av_chipselect -> LEDG:chipselect
	wire          ledg_s1_translator_avalon_anti_slave_0_write;                                                                                     // LEDG_s1_translator:av_write -> LEDG:write_n
	wire   [31:0] ledg_s1_translator_avalon_anti_slave_0_readdata;                                                                                  // LEDG:readdata -> LEDG_s1_translator:av_readdata
	wire   [31:0] ledr_s1_translator_avalon_anti_slave_0_writedata;                                                                                 // LEDR_s1_translator:av_writedata -> LEDR:writedata
	wire    [1:0] ledr_s1_translator_avalon_anti_slave_0_address;                                                                                   // LEDR_s1_translator:av_address -> LEDR:address
	wire          ledr_s1_translator_avalon_anti_slave_0_chipselect;                                                                                // LEDR_s1_translator:av_chipselect -> LEDR:chipselect
	wire          ledr_s1_translator_avalon_anti_slave_0_write;                                                                                     // LEDR_s1_translator:av_write -> LEDR:write_n
	wire   [31:0] ledr_s1_translator_avalon_anti_slave_0_readdata;                                                                                  // LEDR:readdata -> LEDR_s1_translator:av_readdata
	wire    [1:0] switches_s1_translator_avalon_anti_slave_0_address;                                                                               // switches_s1_translator:av_address -> switches:address
	wire   [31:0] switches_s1_translator_avalon_anti_slave_0_readdata;                                                                              // switches:readdata -> switches_s1_translator:av_readdata
	wire    [1:0] key_s1_translator_avalon_anti_slave_0_address;                                                                                    // key_s1_translator:av_address -> key:address
	wire   [31:0] key_s1_translator_avalon_anti_slave_0_readdata;                                                                                   // key:readdata -> key_s1_translator:av_readdata
	wire   [15:0] sdcard_timer_s1_translator_avalon_anti_slave_0_writedata;                                                                         // sdcard_timer_s1_translator:av_writedata -> sdcard_timer:writedata
	wire    [2:0] sdcard_timer_s1_translator_avalon_anti_slave_0_address;                                                                           // sdcard_timer_s1_translator:av_address -> sdcard_timer:address
	wire          sdcard_timer_s1_translator_avalon_anti_slave_0_chipselect;                                                                        // sdcard_timer_s1_translator:av_chipselect -> sdcard_timer:chipselect
	wire          sdcard_timer_s1_translator_avalon_anti_slave_0_write;                                                                             // sdcard_timer_s1_translator:av_write -> sdcard_timer:write_n
	wire   [15:0] sdcard_timer_s1_translator_avalon_anti_slave_0_readdata;                                                                          // sdcard_timer:readdata -> sdcard_timer_s1_translator:av_readdata
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_waitrequest;                              // Altera_UP_SD_Card_Avalon_Interface_0:o_avalon_waitrequest -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:av_waitrequest
	wire   [31:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_writedata;                                // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:av_writedata -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_writedata
	wire    [7:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_address;                                  // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:av_address -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_address
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_chipselect;                               // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:av_chipselect -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_chip_select
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_write;                                    // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:av_write -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_write
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_read;                                     // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:av_read -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_read
	wire   [31:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_readdata;                                 // Altera_UP_SD_Card_Avalon_Interface_0:o_avalon_readdata -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:av_readdata
	wire    [3:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_byteenable;                               // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:av_byteenable -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_byteenable
	wire          ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_waitrequest;                                                                // ps2_0:waitrequest -> ps2_0_avalon_ps2_slave_translator:av_waitrequest
	wire   [31:0] ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_writedata;                                                                  // ps2_0_avalon_ps2_slave_translator:av_writedata -> ps2_0:writedata
	wire    [0:0] ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_address;                                                                    // ps2_0_avalon_ps2_slave_translator:av_address -> ps2_0:address
	wire          ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_chipselect;                                                                 // ps2_0_avalon_ps2_slave_translator:av_chipselect -> ps2_0:chipselect
	wire          ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_write;                                                                      // ps2_0_avalon_ps2_slave_translator:av_write -> ps2_0:write
	wire          ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_read;                                                                       // ps2_0_avalon_ps2_slave_translator:av_read -> ps2_0:read
	wire   [31:0] ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_readdata;                                                                   // ps2_0:readdata -> ps2_0_avalon_ps2_slave_translator:av_readdata
	wire    [3:0] ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_byteenable;                                                                 // ps2_0_avalon_ps2_slave_translator:av_byteenable -> ps2_0:byteenable
	wire   [31:0] audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_writedata;                                                              // audio_0_avalon_audio_slave_translator:av_writedata -> audio_0:writedata
	wire    [1:0] audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_address;                                                                // audio_0_avalon_audio_slave_translator:av_address -> audio_0:address
	wire          audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_chipselect;                                                             // audio_0_avalon_audio_slave_translator:av_chipselect -> audio_0:chipselect
	wire          audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_write;                                                                  // audio_0_avalon_audio_slave_translator:av_write -> audio_0:write
	wire          audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_read;                                                                   // audio_0_avalon_audio_slave_translator:av_read -> audio_0:read
	wire   [31:0] audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_readdata;                                                               // audio_0:readdata -> audio_0_avalon_audio_slave_translator:av_readdata
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_waitrequest;                                                      // character_lcd_0:waitrequest -> character_lcd_0_avalon_lcd_slave_translator:av_waitrequest
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_writedata;                                                        // character_lcd_0_avalon_lcd_slave_translator:av_writedata -> character_lcd_0:writedata
	wire    [0:0] character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_address;                                                          // character_lcd_0_avalon_lcd_slave_translator:av_address -> character_lcd_0:address
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_chipselect;                                                       // character_lcd_0_avalon_lcd_slave_translator:av_chipselect -> character_lcd_0:chipselect
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_write;                                                            // character_lcd_0_avalon_lcd_slave_translator:av_write -> character_lcd_0:write
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_read;                                                             // character_lcd_0_avalon_lcd_slave_translator:av_read -> character_lcd_0:read
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_readdata;                                                         // character_lcd_0:readdata -> character_lcd_0_avalon_lcd_slave_translator:av_readdata
	wire          jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                                                // JTAG:av_waitrequest -> JTAG_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                                                  // JTAG_avalon_jtag_slave_translator:av_writedata -> JTAG:av_writedata
	wire    [0:0] jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                                                    // JTAG_avalon_jtag_slave_translator:av_address -> JTAG:av_address
	wire          jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                                                 // JTAG_avalon_jtag_slave_translator:av_chipselect -> JTAG:av_chipselect
	wire          jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                                                      // JTAG_avalon_jtag_slave_translator:av_write -> JTAG:av_write_n
	wire          jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                                                       // JTAG_avalon_jtag_slave_translator:av_read -> JTAG:av_read_n
	wire   [31:0] jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                                                   // JTAG:av_readdata -> JTAG_avalon_jtag_slave_translator:av_readdata
	wire   [31:0] video_pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_writedata;                                             // video_pixel_buffer_dma_avalon_control_slave_translator:av_writedata -> video_pixel_buffer_dma:slave_writedata
	wire    [1:0] video_pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_address;                                               // video_pixel_buffer_dma_avalon_control_slave_translator:av_address -> video_pixel_buffer_dma:slave_address
	wire          video_pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_write;                                                 // video_pixel_buffer_dma_avalon_control_slave_translator:av_write -> video_pixel_buffer_dma:slave_write
	wire          video_pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_read;                                                  // video_pixel_buffer_dma_avalon_control_slave_translator:av_read -> video_pixel_buffer_dma:slave_read
	wire   [31:0] video_pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_readdata;                                              // video_pixel_buffer_dma:slave_readdata -> video_pixel_buffer_dma_avalon_control_slave_translator:av_readdata
	wire    [3:0] video_pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_byteenable;                                            // video_pixel_buffer_dma_avalon_control_slave_translator:av_byteenable -> video_pixel_buffer_dma:slave_byteenable
	wire   [31:0] video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_anti_slave_0_writedata;                             // video_character_buffer_with_dma_0_avalon_char_control_slave_translator:av_writedata -> video_character_buffer_with_dma_0:ctrl_writedata
	wire    [0:0] video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_anti_slave_0_address;                               // video_character_buffer_with_dma_0_avalon_char_control_slave_translator:av_address -> video_character_buffer_with_dma_0:ctrl_address
	wire          video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_anti_slave_0_chipselect;                            // video_character_buffer_with_dma_0_avalon_char_control_slave_translator:av_chipselect -> video_character_buffer_with_dma_0:ctrl_chipselect
	wire          video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_anti_slave_0_write;                                 // video_character_buffer_with_dma_0_avalon_char_control_slave_translator:av_write -> video_character_buffer_with_dma_0:ctrl_write
	wire          video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_anti_slave_0_read;                                  // video_character_buffer_with_dma_0_avalon_char_control_slave_translator:av_read -> video_character_buffer_with_dma_0:ctrl_read
	wire   [31:0] video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_anti_slave_0_readdata;                              // video_character_buffer_with_dma_0:ctrl_readdata -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator:av_readdata
	wire    [3:0] video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_anti_slave_0_byteenable;                            // video_character_buffer_with_dma_0_avalon_char_control_slave_translator:av_byteenable -> video_character_buffer_with_dma_0:ctrl_byteenable
	wire          video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_anti_slave_0_waitrequest;                            // video_character_buffer_with_dma_0:buf_waitrequest -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator:av_waitrequest
	wire    [7:0] video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_anti_slave_0_writedata;                              // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator:av_writedata -> video_character_buffer_with_dma_0:buf_writedata
	wire   [12:0] video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_anti_slave_0_address;                                // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator:av_address -> video_character_buffer_with_dma_0:buf_address
	wire          video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_anti_slave_0_chipselect;                             // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator:av_chipselect -> video_character_buffer_with_dma_0:buf_chipselect
	wire          video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_anti_slave_0_write;                                  // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator:av_write -> video_character_buffer_with_dma_0:buf_write
	wire          video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_anti_slave_0_read;                                   // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator:av_read -> video_character_buffer_with_dma_0:buf_read
	wire    [7:0] video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_anti_slave_0_readdata;                               // video_character_buffer_with_dma_0:buf_readdata -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator:av_readdata
	wire    [0:0] video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_anti_slave_0_byteenable;                             // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator:av_byteenable -> video_character_buffer_with_dma_0:buf_byteenable
	wire   [15:0] sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_writedata;                                                                // sram_0_avalon_sram_slave_translator:av_writedata -> sram_0:writedata
	wire   [17:0] sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_address;                                                                  // sram_0_avalon_sram_slave_translator:av_address -> sram_0:address
	wire          sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_write;                                                                    // sram_0_avalon_sram_slave_translator:av_write -> sram_0:write
	wire          sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_read;                                                                     // sram_0_avalon_sram_slave_translator:av_read -> sram_0:read
	wire   [15:0] sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_readdata;                                                                 // sram_0:readdata -> sram_0_avalon_sram_slave_translator:av_readdata
	wire          sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid;                                                            // sram_0:readdatavalid -> sram_0_avalon_sram_slave_translator:av_readdatavalid
	wire    [1:0] sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable;                                                               // sram_0_avalon_sram_slave_translator:av_byteenable -> sram_0:byteenable
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest;                                       // audio_and_video_config_0:waitrequest -> audio_and_video_config_0_avalon_av_config_slave_translator:av_waitrequest
	wire   [31:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata;                                         // audio_and_video_config_0_avalon_av_config_slave_translator:av_writedata -> audio_and_video_config_0:writedata
	wire    [1:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_address;                                           // audio_and_video_config_0_avalon_av_config_slave_translator:av_address -> audio_and_video_config_0:address
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_write;                                             // audio_and_video_config_0_avalon_av_config_slave_translator:av_write -> audio_and_video_config_0:write
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_read;                                              // audio_and_video_config_0_avalon_av_config_slave_translator:av_read -> audio_and_video_config_0:read
	wire   [31:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata;                                          // audio_and_video_config_0:readdata -> audio_and_video_config_0_avalon_av_config_slave_translator:av_readdata
	wire    [3:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable;                                        // audio_and_video_config_0_avalon_av_config_slave_translator:av_byteenable -> audio_and_video_config_0:byteenable
	wire   [15:0] usb_0_avalon_usb_slave_translator_avalon_anti_slave_0_writedata;                                                                  // usb_0_avalon_usb_slave_translator:av_writedata -> usb_0:writedata
	wire    [1:0] usb_0_avalon_usb_slave_translator_avalon_anti_slave_0_address;                                                                    // usb_0_avalon_usb_slave_translator:av_address -> usb_0:address
	wire          usb_0_avalon_usb_slave_translator_avalon_anti_slave_0_chipselect;                                                                 // usb_0_avalon_usb_slave_translator:av_chipselect -> usb_0:chipselect
	wire          usb_0_avalon_usb_slave_translator_avalon_anti_slave_0_write;                                                                      // usb_0_avalon_usb_slave_translator:av_write -> usb_0:write
	wire          usb_0_avalon_usb_slave_translator_avalon_anti_slave_0_read;                                                                       // usb_0_avalon_usb_slave_translator:av_read -> usb_0:read
	wire   [15:0] usb_0_avalon_usb_slave_translator_avalon_anti_slave_0_readdata;                                                                   // usb_0:readdata -> usb_0_avalon_usb_slave_translator:av_readdata
	wire          nios2_system_instruction_master_translator_avalon_universal_master_0_waitrequest;                                                 // nios2_system_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_system_instruction_master_translator:uav_waitrequest
	wire    [2:0] nios2_system_instruction_master_translator_avalon_universal_master_0_burstcount;                                                  // nios2_system_instruction_master_translator:uav_burstcount -> nios2_system_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_system_instruction_master_translator_avalon_universal_master_0_writedata;                                                   // nios2_system_instruction_master_translator:uav_writedata -> nios2_system_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] nios2_system_instruction_master_translator_avalon_universal_master_0_address;                                                     // nios2_system_instruction_master_translator:uav_address -> nios2_system_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_system_instruction_master_translator_avalon_universal_master_0_lock;                                                        // nios2_system_instruction_master_translator:uav_lock -> nios2_system_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_system_instruction_master_translator_avalon_universal_master_0_write;                                                       // nios2_system_instruction_master_translator:uav_write -> nios2_system_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_system_instruction_master_translator_avalon_universal_master_0_read;                                                        // nios2_system_instruction_master_translator:uav_read -> nios2_system_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_system_instruction_master_translator_avalon_universal_master_0_readdata;                                                    // nios2_system_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_system_instruction_master_translator:uav_readdata
	wire          nios2_system_instruction_master_translator_avalon_universal_master_0_debugaccess;                                                 // nios2_system_instruction_master_translator:uav_debugaccess -> nios2_system_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_system_instruction_master_translator_avalon_universal_master_0_byteenable;                                                  // nios2_system_instruction_master_translator:uav_byteenable -> nios2_system_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_system_instruction_master_translator_avalon_universal_master_0_readdatavalid;                                               // nios2_system_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_system_instruction_master_translator:uav_readdatavalid
	wire          nios2_system_data_master_translator_avalon_universal_master_0_waitrequest;                                                        // nios2_system_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_system_data_master_translator:uav_waitrequest
	wire    [2:0] nios2_system_data_master_translator_avalon_universal_master_0_burstcount;                                                         // nios2_system_data_master_translator:uav_burstcount -> nios2_system_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_system_data_master_translator_avalon_universal_master_0_writedata;                                                          // nios2_system_data_master_translator:uav_writedata -> nios2_system_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] nios2_system_data_master_translator_avalon_universal_master_0_address;                                                            // nios2_system_data_master_translator:uav_address -> nios2_system_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_system_data_master_translator_avalon_universal_master_0_lock;                                                               // nios2_system_data_master_translator:uav_lock -> nios2_system_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_system_data_master_translator_avalon_universal_master_0_write;                                                              // nios2_system_data_master_translator:uav_write -> nios2_system_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_system_data_master_translator_avalon_universal_master_0_read;                                                               // nios2_system_data_master_translator:uav_read -> nios2_system_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_system_data_master_translator_avalon_universal_master_0_readdata;                                                           // nios2_system_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_system_data_master_translator:uav_readdata
	wire          nios2_system_data_master_translator_avalon_universal_master_0_debugaccess;                                                        // nios2_system_data_master_translator:uav_debugaccess -> nios2_system_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_system_data_master_translator_avalon_universal_master_0_byteenable;                                                         // nios2_system_data_master_translator:uav_byteenable -> nios2_system_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_system_data_master_translator_avalon_universal_master_0_readdatavalid;                                                      // nios2_system_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_system_data_master_translator:uav_readdatavalid
	wire          video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest;                                  // video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_waitrequest -> video_pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_waitrequest
	wire    [1:0] video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount;                                   // video_pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_burstcount -> video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [15:0] video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata;                                    // video_pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_writedata -> video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_address;                                      // video_pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_address -> video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_address
	wire          video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock;                                         // video_pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_lock -> video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_lock
	wire          video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_write;                                        // video_pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_write -> video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_write
	wire          video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_read;                                         // video_pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_read -> video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_read
	wire   [15:0] video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata;                                     // video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_readdata -> video_pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_readdata
	wire          video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess;                                  // video_pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_debugaccess -> video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [1:0] video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable;                                   // video_pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_byteenable -> video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid;                                // video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> video_pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_readdatavalid
	wire          nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                          // nios2_system_jtag_debug_module_translator:uav_waitrequest -> nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                                           // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_system_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                                            // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_system_jtag_debug_module_translator:uav_writedata
	wire   [31:0] nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                                              // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_system_jtag_debug_module_translator:uav_address
	wire          nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                                                // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_system_jtag_debug_module_translator:uav_write
	wire          nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                                                 // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_system_jtag_debug_module_translator:uav_lock
	wire          nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                                                 // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_system_jtag_debug_module_translator:uav_read
	wire   [31:0] nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                                             // nios2_system_jtag_debug_module_translator:uav_readdata -> nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                        // nios2_system_jtag_debug_module_translator:uav_readdatavalid -> nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                          // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_system_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                                           // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_system_jtag_debug_module_translator:uav_byteenable
	wire          nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                   // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                                         // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                 // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                                          // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                                         // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                      // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                              // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                       // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                      // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                    // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                     // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                    // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          onchip_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                               // onchip_s1_translator:uav_waitrequest -> onchip_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] onchip_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                                // onchip_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_s1_translator:uav_burstcount
	wire   [31:0] onchip_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                                 // onchip_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_s1_translator:uav_writedata
	wire   [31:0] onchip_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                                   // onchip_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_s1_translator:uav_address
	wire          onchip_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                                     // onchip_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_s1_translator:uav_write
	wire          onchip_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                                      // onchip_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_s1_translator:uav_lock
	wire          onchip_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                                      // onchip_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_s1_translator:uav_read
	wire   [31:0] onchip_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                                  // onchip_s1_translator:uav_readdata -> onchip_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          onchip_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                             // onchip_s1_translator:uav_readdatavalid -> onchip_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          onchip_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                               // onchip_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_s1_translator:uav_debugaccess
	wire    [3:0] onchip_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                                // onchip_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_s1_translator:uav_byteenable
	wire          onchip_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                                        // onchip_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          onchip_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                              // onchip_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          onchip_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                                      // onchip_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] onchip_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                               // onchip_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          onchip_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                              // onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                                     // onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                           // onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                                   // onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                            // onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                           // onchip_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          onchip_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                                         // onchip_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] onchip_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                          // onchip_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          onchip_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                                         // onchip_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                                // sdram_s1_translator:uav_waitrequest -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                                 // sdram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_s1_translator:uav_burstcount
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                                  // sdram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_s1_translator:uav_writedata
	wire   [31:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                                    // sdram_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_s1_translator:uav_address
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                                      // sdram_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_s1_translator:uav_write
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                                       // sdram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_s1_translator:uav_lock
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                                       // sdram_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_s1_translator:uav_read
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                                   // sdram_s1_translator:uav_readdata -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                              // sdram_s1_translator:uav_readdatavalid -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                                // sdram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_s1_translator:uav_debugaccess
	wire    [1:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                                 // sdram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_s1_translator:uav_byteenable
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                                         // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                               // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                                       // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [91:0] sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                                // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                               // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                                      // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                            // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                                    // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [91:0] sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                             // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                            // sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                                          // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [17:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                           // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                                          // sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                                          // sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [17:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                                           // sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                                          // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                                 // LEDG_s1_translator:uav_waitrequest -> LEDG_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ledg_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                                  // LEDG_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> LEDG_s1_translator:uav_burstcount
	wire   [31:0] ledg_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                                   // LEDG_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> LEDG_s1_translator:uav_writedata
	wire   [31:0] ledg_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                                     // LEDG_s1_translator_avalon_universal_slave_0_agent:m0_address -> LEDG_s1_translator:uav_address
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                                       // LEDG_s1_translator_avalon_universal_slave_0_agent:m0_write -> LEDG_s1_translator:uav_write
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                                        // LEDG_s1_translator_avalon_universal_slave_0_agent:m0_lock -> LEDG_s1_translator:uav_lock
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                                        // LEDG_s1_translator_avalon_universal_slave_0_agent:m0_read -> LEDG_s1_translator:uav_read
	wire   [31:0] ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                                    // LEDG_s1_translator:uav_readdata -> LEDG_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                               // LEDG_s1_translator:uav_readdatavalid -> LEDG_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                                 // LEDG_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> LEDG_s1_translator:uav_debugaccess
	wire    [3:0] ledg_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                                  // LEDG_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> LEDG_s1_translator:uav_byteenable
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                                          // LEDG_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                                // LEDG_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                                        // LEDG_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                                 // LEDG_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                                // LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> LEDG_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                                       // LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> LEDG_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                             // LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> LEDG_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                                     // LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> LEDG_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                              // LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> LEDG_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                             // LEDG_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                                           // LEDG_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> LEDG_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                            // LEDG_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> LEDG_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                                           // LEDG_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> LEDG_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                                 // LEDR_s1_translator:uav_waitrequest -> LEDR_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                                  // LEDR_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> LEDR_s1_translator:uav_burstcount
	wire   [31:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                                   // LEDR_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> LEDR_s1_translator:uav_writedata
	wire   [31:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                                     // LEDR_s1_translator_avalon_universal_slave_0_agent:m0_address -> LEDR_s1_translator:uav_address
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                                       // LEDR_s1_translator_avalon_universal_slave_0_agent:m0_write -> LEDR_s1_translator:uav_write
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                                        // LEDR_s1_translator_avalon_universal_slave_0_agent:m0_lock -> LEDR_s1_translator:uav_lock
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                                        // LEDR_s1_translator_avalon_universal_slave_0_agent:m0_read -> LEDR_s1_translator:uav_read
	wire   [31:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                                    // LEDR_s1_translator:uav_readdata -> LEDR_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                               // LEDR_s1_translator:uav_readdatavalid -> LEDR_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                                 // LEDR_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> LEDR_s1_translator:uav_debugaccess
	wire    [3:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                                  // LEDR_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> LEDR_s1_translator:uav_byteenable
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                                          // LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                                // LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                                        // LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                                 // LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                                // LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                                       // LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                             // LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                                     // LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                              // LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                             // LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                                           // LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                            // LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                                           // LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          switches_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                             // switches_s1_translator:uav_waitrequest -> switches_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                              // switches_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> switches_s1_translator:uav_burstcount
	wire   [31:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                               // switches_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> switches_s1_translator:uav_writedata
	wire   [31:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                                 // switches_s1_translator_avalon_universal_slave_0_agent:m0_address -> switches_s1_translator:uav_address
	wire          switches_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                                   // switches_s1_translator_avalon_universal_slave_0_agent:m0_write -> switches_s1_translator:uav_write
	wire          switches_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                                    // switches_s1_translator_avalon_universal_slave_0_agent:m0_lock -> switches_s1_translator:uav_lock
	wire          switches_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                                    // switches_s1_translator_avalon_universal_slave_0_agent:m0_read -> switches_s1_translator:uav_read
	wire   [31:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                                // switches_s1_translator:uav_readdata -> switches_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          switches_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                           // switches_s1_translator:uav_readdatavalid -> switches_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          switches_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                             // switches_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> switches_s1_translator:uav_debugaccess
	wire    [3:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                              // switches_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> switches_s1_translator:uav_byteenable
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                                      // switches_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                            // switches_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                                    // switches_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] switches_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                             // switches_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                            // switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> switches_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                                   // switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                         // switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                                 // switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                          // switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                         // switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                                       // switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                        // switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                                       // switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          key_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                                  // key_s1_translator:uav_waitrequest -> key_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] key_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                                   // key_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> key_s1_translator:uav_burstcount
	wire   [31:0] key_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                                    // key_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> key_s1_translator:uav_writedata
	wire   [31:0] key_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                                      // key_s1_translator_avalon_universal_slave_0_agent:m0_address -> key_s1_translator:uav_address
	wire          key_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                                        // key_s1_translator_avalon_universal_slave_0_agent:m0_write -> key_s1_translator:uav_write
	wire          key_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                                         // key_s1_translator_avalon_universal_slave_0_agent:m0_lock -> key_s1_translator:uav_lock
	wire          key_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                                         // key_s1_translator_avalon_universal_slave_0_agent:m0_read -> key_s1_translator:uav_read
	wire   [31:0] key_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                                     // key_s1_translator:uav_readdata -> key_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          key_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                                // key_s1_translator:uav_readdatavalid -> key_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          key_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                                  // key_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> key_s1_translator:uav_debugaccess
	wire    [3:0] key_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                                   // key_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> key_s1_translator:uav_byteenable
	wire          key_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                                           // key_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          key_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                                 // key_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          key_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                                         // key_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] key_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                                  // key_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          key_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                                 // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> key_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                                        // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> key_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                              // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> key_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                                      // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> key_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                               // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> key_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                              // key_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                                            // key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                             // key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                                            // key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                         // sdcard_timer_s1_translator:uav_waitrequest -> sdcard_timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                          // sdcard_timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdcard_timer_s1_translator:uav_burstcount
	wire   [31:0] sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                           // sdcard_timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdcard_timer_s1_translator:uav_writedata
	wire   [31:0] sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                             // sdcard_timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdcard_timer_s1_translator:uav_address
	wire          sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                               // sdcard_timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdcard_timer_s1_translator:uav_write
	wire          sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                                // sdcard_timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdcard_timer_s1_translator:uav_lock
	wire          sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                                // sdcard_timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdcard_timer_s1_translator:uav_read
	wire   [31:0] sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                            // sdcard_timer_s1_translator:uav_readdata -> sdcard_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                       // sdcard_timer_s1_translator:uav_readdatavalid -> sdcard_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                         // sdcard_timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdcard_timer_s1_translator:uav_debugaccess
	wire    [3:0] sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                          // sdcard_timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdcard_timer_s1_translator:uav_byteenable
	wire          sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                                  // sdcard_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                        // sdcard_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                                // sdcard_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                         // sdcard_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                        // sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdcard_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                               // sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdcard_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                     // sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdcard_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                             // sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdcard_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                      // sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdcard_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                     // sdcard_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                                   // sdcard_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdcard_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                    // sdcard_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdcard_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                                   // sdcard_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdcard_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_waitrequest -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                 // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_burstcount
	wire   [31:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                  // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_writedata
	wire   [31:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_address;                    // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_address -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_address
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_write;                      // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_write -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_write
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_lock;                       // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_lock
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_read;                       // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_read -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_read
	wire   [31:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                   // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_readdata -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;              // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_readdatavalid -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_debugaccess
	wire    [3:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                 // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_byteenable
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;         // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;               // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;       // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;               // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;      // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;            // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;    // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;             // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;            // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;          // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;           // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;          // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                  // ps2_0_avalon_ps2_slave_translator:uav_waitrequest -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                   // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> ps2_0_avalon_ps2_slave_translator:uav_burstcount
	wire   [31:0] ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                                    // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> ps2_0_avalon_ps2_slave_translator:uav_writedata
	wire   [31:0] ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_address;                                                      // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_address -> ps2_0_avalon_ps2_slave_translator:uav_address
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_write;                                                        // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_write -> ps2_0_avalon_ps2_slave_translator:uav_write
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                                         // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_lock -> ps2_0_avalon_ps2_slave_translator:uav_lock
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_read;                                                         // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_read -> ps2_0_avalon_ps2_slave_translator:uav_read
	wire   [31:0] ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                                     // ps2_0_avalon_ps2_slave_translator:uav_readdata -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                // ps2_0_avalon_ps2_slave_translator:uav_readdatavalid -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                  // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ps2_0_avalon_ps2_slave_translator:uav_debugaccess
	wire    [3:0] ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                   // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> ps2_0_avalon_ps2_slave_translator:uav_byteenable
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                           // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                 // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                         // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                                  // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                 // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                        // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                              // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                      // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                               // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                              // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                            // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                             // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                            // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                              // audio_0_avalon_audio_slave_translator:uav_waitrequest -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                               // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> audio_0_avalon_audio_slave_translator:uav_burstcount
	wire   [31:0] audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                                // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> audio_0_avalon_audio_slave_translator:uav_writedata
	wire   [31:0] audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_address;                                                  // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_address -> audio_0_avalon_audio_slave_translator:uav_address
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_write;                                                    // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_write -> audio_0_avalon_audio_slave_translator:uav_write
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                                     // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_lock -> audio_0_avalon_audio_slave_translator:uav_lock
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_read;                                                     // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_read -> audio_0_avalon_audio_slave_translator:uav_read
	wire   [31:0] audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                                 // audio_0_avalon_audio_slave_translator:uav_readdata -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                            // audio_0_avalon_audio_slave_translator:uav_readdatavalid -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                              // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> audio_0_avalon_audio_slave_translator:uav_debugaccess
	wire    [3:0] audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                               // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> audio_0_avalon_audio_slave_translator:uav_byteenable
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                       // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                             // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                     // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                              // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                             // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                    // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                          // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                  // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                           // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                          // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                        // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                         // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                        // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                        // character_lcd_0_avalon_lcd_slave_translator:uav_waitrequest -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [0:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                         // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> character_lcd_0_avalon_lcd_slave_translator:uav_burstcount
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                          // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> character_lcd_0_avalon_lcd_slave_translator:uav_writedata
	wire   [31:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_address;                                            // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_address -> character_lcd_0_avalon_lcd_slave_translator:uav_address
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_write;                                              // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_write -> character_lcd_0_avalon_lcd_slave_translator:uav_write
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                               // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_lock -> character_lcd_0_avalon_lcd_slave_translator:uav_lock
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_read;                                               // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_read -> character_lcd_0_avalon_lcd_slave_translator:uav_read
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                           // character_lcd_0_avalon_lcd_slave_translator:uav_readdata -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                      // character_lcd_0_avalon_lcd_slave_translator:uav_readdatavalid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                        // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> character_lcd_0_avalon_lcd_slave_translator:uav_debugaccess
	wire    [0:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                         // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> character_lcd_0_avalon_lcd_slave_translator:uav_byteenable
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                 // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                       // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                               // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [82:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                        // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                       // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                              // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                    // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                            // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [82:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                     // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                    // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                  // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire    [9:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                   // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                  // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                  // JTAG_avalon_jtag_slave_translator:uav_waitrequest -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                   // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> JTAG_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                                    // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> JTAG_avalon_jtag_slave_translator:uav_writedata
	wire   [31:0] jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                                                      // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> JTAG_avalon_jtag_slave_translator:uav_address
	wire          jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                                                        // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> JTAG_avalon_jtag_slave_translator:uav_write
	wire          jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                                         // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> JTAG_avalon_jtag_slave_translator:uav_lock
	wire          jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                                                         // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> JTAG_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                                     // JTAG_avalon_jtag_slave_translator:uav_readdata -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                // JTAG_avalon_jtag_slave_translator:uav_readdatavalid -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                  // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> JTAG_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                   // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> JTAG_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                           // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                 // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                         // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                                  // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                 // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                        // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                              // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                      // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                               // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                              // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                            // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                             // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                            // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // video_pixel_buffer_dma_avalon_control_slave_translator:uav_waitrequest -> video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> video_pixel_buffer_dma_avalon_control_slave_translator:uav_burstcount
	wire   [31:0] video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                               // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> video_pixel_buffer_dma_avalon_control_slave_translator:uav_writedata
	wire   [31:0] video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                                 // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> video_pixel_buffer_dma_avalon_control_slave_translator:uav_address
	wire          video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                                   // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> video_pixel_buffer_dma_avalon_control_slave_translator:uav_write
	wire          video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                    // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> video_pixel_buffer_dma_avalon_control_slave_translator:uav_lock
	wire          video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                                    // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> video_pixel_buffer_dma_avalon_control_slave_translator:uav_read
	wire   [31:0] video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                // video_pixel_buffer_dma_avalon_control_slave_translator:uav_readdata -> video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // video_pixel_buffer_dma_avalon_control_slave_translator:uav_readdatavalid -> video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> video_pixel_buffer_dma_avalon_control_slave_translator:uav_debugaccess
	wire    [3:0] video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> video_pixel_buffer_dma_avalon_control_slave_translator:uav_byteenable
	wire          video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                             // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // video_character_buffer_with_dma_0_avalon_char_control_slave_translator:uav_waitrequest -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator:uav_burstcount
	wire   [31:0] video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator:uav_writedata
	wire   [31:0] video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator:uav_address
	wire          video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator:uav_write
	wire          video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator:uav_lock
	wire          video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator:uav_read
	wire   [31:0] video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // video_character_buffer_with_dma_0_avalon_char_control_slave_translator:uav_readdata -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // video_character_buffer_with_dma_0_avalon_char_control_slave_translator:uav_readdatavalid -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator:uav_debugaccess
	wire    [3:0] video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator:uav_byteenable
	wire          video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator:uav_waitrequest -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [0:0] video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;               // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator:uav_burstcount
	wire    [7:0] video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator:uav_writedata
	wire   [31:0] video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_address;                  // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_address -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator:uav_address
	wire          video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_write;                    // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_write -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator:uav_write
	wire          video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_lock;                     // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_lock -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator:uav_lock
	wire          video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_read;                     // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_read -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator:uav_read
	wire    [7:0] video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                 // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator:uav_readdata -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator:uav_readdatavalid -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator:uav_debugaccess
	wire    [0:0] video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;               // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator:uav_byteenable
	wire          video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;             // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [82:0] video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_data;              // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;             // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [82:0] video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire    [9:0] video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                // sram_0_avalon_sram_slave_translator:uav_waitrequest -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                 // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sram_0_avalon_sram_slave_translator:uav_burstcount
	wire   [15:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                                  // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sram_0_avalon_sram_slave_translator:uav_writedata
	wire   [31:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address;                                                    // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_address -> sram_0_avalon_sram_slave_translator:uav_address
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write;                                                      // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_write -> sram_0_avalon_sram_slave_translator:uav_write
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                                       // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sram_0_avalon_sram_slave_translator:uav_lock
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read;                                                       // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_read -> sram_0_avalon_sram_slave_translator:uav_read
	wire   [15:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                                   // sram_0_avalon_sram_slave_translator:uav_readdata -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                              // sram_0_avalon_sram_slave_translator:uav_readdatavalid -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sram_0_avalon_sram_slave_translator:uav_debugaccess
	wire    [1:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                 // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sram_0_avalon_sram_slave_translator:uav_byteenable
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                         // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                               // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                       // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [91:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                                // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                               // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                      // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                            // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                    // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [91:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                             // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                            // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                          // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [17:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                           // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                          // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                          // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [17:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                           // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                          // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // audio_and_video_config_0_avalon_av_config_slave_translator:uav_waitrequest -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_burstcount
	wire   [31:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                           // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_writedata
	wire   [31:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address;                             // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_address -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_address
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write;                               // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_write -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_write
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_lock -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_lock
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read;                                // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_read -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_read
	wire   [31:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                            // audio_and_video_config_0_avalon_av_config_slave_translator:uav_readdata -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // audio_and_video_config_0_avalon_av_config_slave_translator:uav_readdatavalid -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_debugaccess
	wire    [3:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> audio_and_video_config_0_avalon_av_config_slave_translator:uav_byteenable
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                         // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                  // usb_0_avalon_usb_slave_translator:uav_waitrequest -> usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                   // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> usb_0_avalon_usb_slave_translator:uav_burstcount
	wire   [31:0] usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                                    // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> usb_0_avalon_usb_slave_translator:uav_writedata
	wire   [31:0] usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_address;                                                      // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:m0_address -> usb_0_avalon_usb_slave_translator:uav_address
	wire          usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_write;                                                        // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:m0_write -> usb_0_avalon_usb_slave_translator:uav_write
	wire          usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                                         // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:m0_lock -> usb_0_avalon_usb_slave_translator:uav_lock
	wire          usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_read;                                                         // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:m0_read -> usb_0_avalon_usb_slave_translator:uav_read
	wire   [31:0] usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                                     // usb_0_avalon_usb_slave_translator:uav_readdata -> usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                // usb_0_avalon_usb_slave_translator:uav_readdatavalid -> usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                  // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> usb_0_avalon_usb_slave_translator:uav_debugaccess
	wire    [3:0] usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                   // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> usb_0_avalon_usb_slave_translator:uav_byteenable
	wire          usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                           // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                 // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                         // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                                  // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                 // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                        // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                              // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                      // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                               // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                              // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                            // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                             // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                            // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          nios2_system_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                                        // nios2_system_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          nios2_system_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                                              // nios2_system_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          nios2_system_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                                      // nios2_system_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [108:0] nios2_system_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                                               // nios2_system_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          nios2_system_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                                              // addr_router:sink_ready -> nios2_system_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_system_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                                               // nios2_system_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          nios2_system_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                                     // nios2_system_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          nios2_system_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                                             // nios2_system_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [108:0] nios2_system_data_master_translator_avalon_universal_master_0_agent_cp_data;                                                      // nios2_system_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          nios2_system_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                                     // addr_router_001:sink_ready -> nios2_system_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                         // video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid;                               // video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                       // video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire   [90:0] video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data;                                // video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready;                               // addr_router_002:sink_ready -> video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                          // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                                                // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                        // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [108:0] nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                                                 // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                                                // id_router:sink_ready -> nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          onchip_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                               // onchip_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          onchip_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                                     // onchip_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          onchip_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                             // onchip_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [108:0] onchip_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                                      // onchip_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          onchip_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                                     // id_router_001:sink_ready -> onchip_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                                // sdram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                                      // sdram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                              // sdram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire   [90:0] sdram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                                       // sdram_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                                      // id_router_002:sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                                 // LEDG_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                                       // LEDG_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                               // LEDG_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [108:0] ledg_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                                        // LEDG_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          ledg_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                                       // id_router_003:sink_ready -> LEDG_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                                 // LEDR_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                                       // LEDR_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                               // LEDR_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [108:0] ledr_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                                        // LEDR_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                                       // id_router_004:sink_ready -> LEDR_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                             // switches_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                                   // switches_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                           // switches_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [108:0] switches_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                                    // switches_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                                   // id_router_005:sink_ready -> switches_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          key_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                                  // key_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          key_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                                        // key_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          key_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                                // key_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [108:0] key_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                                         // key_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          key_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                                        // id_router_006:sink_ready -> key_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                         // sdcard_timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                               // sdcard_timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                       // sdcard_timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [108:0] sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                                // sdcard_timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                               // id_router_007:sink_ready -> sdcard_timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_valid;                      // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;              // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [108:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_data;                       // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_ready;                      // id_router_008:sink_ready -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                  // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                                        // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [108:0] ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_data;                                                         // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                                        // id_router_009:sink_ready -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                              // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                                    // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                            // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [108:0] audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_data;                                                     // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                                    // id_router_010:sink_ready -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                        // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                              // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                      // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire   [81:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_data;                                               // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                              // id_router_011:sink_ready -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                  // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                                        // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [108:0] jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                                                         // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                                        // id_router_012:sink_ready -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                   // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [108:0] video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                                    // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_013:sink_ready -> video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire          video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire          video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire  [108:0] video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire          video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_014:sink_ready -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire          video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_valid;                    // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire          video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire   [81:0] video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_data;                     // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire          video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_015:sink_ready -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                                      // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                              // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire   [90:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data;                                                       // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire          sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                                      // id_router_016:sink_ready -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid;                               // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire  [108:0] audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data;                                // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire          audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_017:sink_ready -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                  // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	wire          usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                                        // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	wire          usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	wire  [108:0] usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_data;                                                         // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	wire          usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                                        // id_router_018:sink_ready -> usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_src_endofpacket;                                                                                                      // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                                                            // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                                                                    // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [108:0] addr_router_src_data;                                                                                                             // addr_router:src_data -> limiter:cmd_sink_data
	wire   [18:0] addr_router_src_channel;                                                                                                          // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                                                            // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                                                      // limiter:rsp_src_endofpacket -> nios2_system_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                                                            // limiter:rsp_src_valid -> nios2_system_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                                                    // limiter:rsp_src_startofpacket -> nios2_system_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [108:0] limiter_rsp_src_data;                                                                                                             // limiter:rsp_src_data -> nios2_system_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [18:0] limiter_rsp_src_channel;                                                                                                          // limiter:rsp_src_channel -> nios2_system_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                                                            // nios2_system_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          addr_router_001_src_endofpacket;                                                                                                  // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire          addr_router_001_src_valid;                                                                                                        // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire          addr_router_001_src_startofpacket;                                                                                                // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [108:0] addr_router_001_src_data;                                                                                                         // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire   [18:0] addr_router_001_src_channel;                                                                                                      // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire          addr_router_001_src_ready;                                                                                                        // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire          limiter_001_rsp_src_endofpacket;                                                                                                  // limiter_001:rsp_src_endofpacket -> nios2_system_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_001_rsp_src_valid;                                                                                                        // limiter_001:rsp_src_valid -> nios2_system_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_001_rsp_src_startofpacket;                                                                                                // limiter_001:rsp_src_startofpacket -> nios2_system_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [108:0] limiter_001_rsp_src_data;                                                                                                         // limiter_001:rsp_src_data -> nios2_system_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [18:0] limiter_001_rsp_src_channel;                                                                                                      // limiter_001:rsp_src_channel -> nios2_system_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_001_rsp_src_ready;                                                                                                        // nios2_system_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire          addr_router_002_src_endofpacket;                                                                                                  // addr_router_002:src_endofpacket -> limiter_002:cmd_sink_endofpacket
	wire          addr_router_002_src_valid;                                                                                                        // addr_router_002:src_valid -> limiter_002:cmd_sink_valid
	wire          addr_router_002_src_startofpacket;                                                                                                // addr_router_002:src_startofpacket -> limiter_002:cmd_sink_startofpacket
	wire   [90:0] addr_router_002_src_data;                                                                                                         // addr_router_002:src_data -> limiter_002:cmd_sink_data
	wire   [18:0] addr_router_002_src_channel;                                                                                                      // addr_router_002:src_channel -> limiter_002:cmd_sink_channel
	wire          addr_router_002_src_ready;                                                                                                        // limiter_002:cmd_sink_ready -> addr_router_002:src_ready
	wire          limiter_002_rsp_src_endofpacket;                                                                                                  // limiter_002:rsp_src_endofpacket -> video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_002_rsp_src_valid;                                                                                                        // limiter_002:rsp_src_valid -> video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_002_rsp_src_startofpacket;                                                                                                // limiter_002:rsp_src_startofpacket -> video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [90:0] limiter_002_rsp_src_data;                                                                                                         // limiter_002:rsp_src_data -> video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [18:0] limiter_002_rsp_src_channel;                                                                                                      // limiter_002:rsp_src_channel -> video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_002_rsp_src_ready;                                                                                                        // video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_002:rsp_src_ready
	wire          burst_adapter_source0_endofpacket;                                                                                                // burst_adapter:source0_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                                                      // burst_adapter:source0_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                                              // burst_adapter:source0_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [90:0] burst_adapter_source0_data;                                                                                                       // burst_adapter:source0_data -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                                                      // sdram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [18:0] burst_adapter_source0_channel;                                                                                                    // burst_adapter:source0_channel -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_001_source0_endofpacket;                                                                                            // burst_adapter_001:source0_endofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_001_source0_valid;                                                                                                  // burst_adapter_001:source0_valid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_001_source0_startofpacket;                                                                                          // burst_adapter_001:source0_startofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [81:0] burst_adapter_001_source0_data;                                                                                                   // burst_adapter_001:source0_data -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_001_source0_ready;                                                                                                  // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire   [18:0] burst_adapter_001_source0_channel;                                                                                                // burst_adapter_001:source0_channel -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_002_source0_endofpacket;                                                                                            // burst_adapter_002:source0_endofpacket -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_002_source0_valid;                                                                                                  // burst_adapter_002:source0_valid -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_002_source0_startofpacket;                                                                                          // burst_adapter_002:source0_startofpacket -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [81:0] burst_adapter_002_source0_data;                                                                                                   // burst_adapter_002:source0_data -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_002_source0_ready;                                                                                                  // video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_002:source0_ready
	wire   [18:0] burst_adapter_002_source0_channel;                                                                                                // burst_adapter_002:source0_channel -> video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_003_source0_endofpacket;                                                                                            // burst_adapter_003:source0_endofpacket -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_003_source0_valid;                                                                                                  // burst_adapter_003:source0_valid -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_003_source0_startofpacket;                                                                                          // burst_adapter_003:source0_startofpacket -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [90:0] burst_adapter_003_source0_data;                                                                                                   // burst_adapter_003:source0_data -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_003_source0_ready;                                                                                                  // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_003:source0_ready
	wire   [18:0] burst_adapter_003_source0_channel;                                                                                                // burst_adapter_003:source0_channel -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                                                   // rst_controller:reset_out -> [Altera_UP_SD_Card_Avalon_Interface_0:i_reset_n, Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:reset, Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:reset, Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, JTAG:rst_n, JTAG_avalon_jtag_slave_translator:reset, JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, LEDG:reset_n, LEDG_s1_translator:reset, LEDG_s1_translator_avalon_universal_slave_0_agent:reset, LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, LEDR:reset_n, LEDR_s1_translator:reset, LEDR_s1_translator_avalon_universal_slave_0_agent:reset, LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, addr_router_002:reset, audio_0:reset, audio_0_avalon_audio_slave_translator:reset, audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:reset, audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, audio_and_video_config_0:reset, audio_and_video_config_0_avalon_av_config_slave_translator:reset, audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:reset, audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, burst_adapter:reset, burst_adapter_001:reset, burst_adapter_002:reset, burst_adapter_003:reset, character_lcd_0:reset, character_lcd_0_avalon_lcd_slave_translator:reset, character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:reset, character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_004:reset, cmd_xbar_mux_005:reset, cmd_xbar_mux_006:reset, cmd_xbar_mux_007:reset, cmd_xbar_mux_008:reset, cmd_xbar_mux_009:reset, cmd_xbar_mux_010:reset, cmd_xbar_mux_016:reset, cmd_xbar_mux_018:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, id_router_017:reset, id_router_018:reset, irq_mapper:reset, key:reset_n, key_s1_translator:reset, key_s1_translator_avalon_universal_slave_0_agent:reset, key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, limiter_001:reset, limiter_002:reset, nios2_system:reset_n, nios2_system_data_master_translator:reset, nios2_system_data_master_translator_avalon_universal_master_0_agent:reset, nios2_system_instruction_master_translator:reset, nios2_system_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_system_jtag_debug_module_translator:reset, nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip:reset, onchip_s1_translator:reset, onchip_s1_translator_avalon_universal_slave_0_agent:reset, onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ps2_0:reset, ps2_0_avalon_ps2_slave_translator:reset, ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:reset, ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_018:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rsp_xbar_mux_002:reset, sdcard_timer:reset_n, sdcard_timer_s1_translator:reset, sdcard_timer_s1_translator_avalon_universal_slave_0_agent:reset, sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sdram:reset_n, sdram_s1_translator:reset, sdram_s1_translator_avalon_universal_slave_0_agent:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sram_0:reset, sram_0_avalon_sram_slave_translator:reset, sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:reset, sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, switches:reset_n, switches_s1_translator:reset, switches_s1_translator_avalon_universal_slave_0_agent:reset, switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, usb_0:reset, usb_0_avalon_usb_slave_translator:reset, usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:reset, usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, video_alpha_blender_0:reset, video_character_buffer_with_dma_0:reset, video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator:reset, video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:reset, video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, video_character_buffer_with_dma_0_avalon_char_control_slave_translator:reset, video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:reset, video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, video_dual_clock_buffer_0:reset_stream_in, video_pixel_buffer_dma:reset, video_pixel_buffer_dma_avalon_control_slave_translator:reset, video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:reset, video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, video_pixel_buffer_dma_avalon_pixel_dma_master_translator:reset, video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:reset, video_rgb_resampler_0:reset, video_scaler_0:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset, width_adapter_004:reset, width_adapter_005:reset, width_adapter_006:reset, width_adapter_007:reset, width_adapter_008:reset, width_adapter_009:reset, width_adapter_010:reset, width_adapter_011:reset]
	wire          rst_controller_reset_out_reset_req;                                                                                               // rst_controller:reset_req -> onchip:reset_req
	wire          nios2_system_jtag_debug_module_reset_reset;                                                                                       // nios2_system:jtag_debug_module_resetrequest -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	wire          rst_controller_001_reset_out_reset;                                                                                               // rst_controller_001:reset_out -> clocks:reset
	wire          rst_controller_002_reset_out_reset;                                                                                               // rst_controller_002:reset_out -> [video_dual_clock_buffer_0:reset_stream_out, video_vga_controller_0:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                                                  // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                                                        // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                                                // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [108:0] cmd_xbar_demux_src0_data;                                                                                                         // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [18:0] cmd_xbar_demux_src0_channel;                                                                                                      // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                                                        // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                                                  // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                                                        // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                                                // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [108:0] cmd_xbar_demux_src1_data;                                                                                                         // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [18:0] cmd_xbar_demux_src1_channel;                                                                                                      // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                                                        // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_src3_endofpacket;                                                                                                  // cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire          cmd_xbar_demux_src3_valid;                                                                                                        // cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	wire          cmd_xbar_demux_src3_startofpacket;                                                                                                // cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [108:0] cmd_xbar_demux_src3_data;                                                                                                         // cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	wire   [18:0] cmd_xbar_demux_src3_channel;                                                                                                      // cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	wire          cmd_xbar_demux_src3_ready;                                                                                                        // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	wire          cmd_xbar_demux_src4_endofpacket;                                                                                                  // cmd_xbar_demux:src4_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	wire          cmd_xbar_demux_src4_valid;                                                                                                        // cmd_xbar_demux:src4_valid -> cmd_xbar_mux_004:sink0_valid
	wire          cmd_xbar_demux_src4_startofpacket;                                                                                                // cmd_xbar_demux:src4_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	wire  [108:0] cmd_xbar_demux_src4_data;                                                                                                         // cmd_xbar_demux:src4_data -> cmd_xbar_mux_004:sink0_data
	wire   [18:0] cmd_xbar_demux_src4_channel;                                                                                                      // cmd_xbar_demux:src4_channel -> cmd_xbar_mux_004:sink0_channel
	wire          cmd_xbar_demux_src4_ready;                                                                                                        // cmd_xbar_mux_004:sink0_ready -> cmd_xbar_demux:src4_ready
	wire          cmd_xbar_demux_src5_endofpacket;                                                                                                  // cmd_xbar_demux:src5_endofpacket -> cmd_xbar_mux_005:sink0_endofpacket
	wire          cmd_xbar_demux_src5_valid;                                                                                                        // cmd_xbar_demux:src5_valid -> cmd_xbar_mux_005:sink0_valid
	wire          cmd_xbar_demux_src5_startofpacket;                                                                                                // cmd_xbar_demux:src5_startofpacket -> cmd_xbar_mux_005:sink0_startofpacket
	wire  [108:0] cmd_xbar_demux_src5_data;                                                                                                         // cmd_xbar_demux:src5_data -> cmd_xbar_mux_005:sink0_data
	wire   [18:0] cmd_xbar_demux_src5_channel;                                                                                                      // cmd_xbar_demux:src5_channel -> cmd_xbar_mux_005:sink0_channel
	wire          cmd_xbar_demux_src5_ready;                                                                                                        // cmd_xbar_mux_005:sink0_ready -> cmd_xbar_demux:src5_ready
	wire          cmd_xbar_demux_src6_endofpacket;                                                                                                  // cmd_xbar_demux:src6_endofpacket -> cmd_xbar_mux_006:sink0_endofpacket
	wire          cmd_xbar_demux_src6_valid;                                                                                                        // cmd_xbar_demux:src6_valid -> cmd_xbar_mux_006:sink0_valid
	wire          cmd_xbar_demux_src6_startofpacket;                                                                                                // cmd_xbar_demux:src6_startofpacket -> cmd_xbar_mux_006:sink0_startofpacket
	wire  [108:0] cmd_xbar_demux_src6_data;                                                                                                         // cmd_xbar_demux:src6_data -> cmd_xbar_mux_006:sink0_data
	wire   [18:0] cmd_xbar_demux_src6_channel;                                                                                                      // cmd_xbar_demux:src6_channel -> cmd_xbar_mux_006:sink0_channel
	wire          cmd_xbar_demux_src6_ready;                                                                                                        // cmd_xbar_mux_006:sink0_ready -> cmd_xbar_demux:src6_ready
	wire          cmd_xbar_demux_src7_endofpacket;                                                                                                  // cmd_xbar_demux:src7_endofpacket -> cmd_xbar_mux_007:sink0_endofpacket
	wire          cmd_xbar_demux_src7_valid;                                                                                                        // cmd_xbar_demux:src7_valid -> cmd_xbar_mux_007:sink0_valid
	wire          cmd_xbar_demux_src7_startofpacket;                                                                                                // cmd_xbar_demux:src7_startofpacket -> cmd_xbar_mux_007:sink0_startofpacket
	wire  [108:0] cmd_xbar_demux_src7_data;                                                                                                         // cmd_xbar_demux:src7_data -> cmd_xbar_mux_007:sink0_data
	wire   [18:0] cmd_xbar_demux_src7_channel;                                                                                                      // cmd_xbar_demux:src7_channel -> cmd_xbar_mux_007:sink0_channel
	wire          cmd_xbar_demux_src7_ready;                                                                                                        // cmd_xbar_mux_007:sink0_ready -> cmd_xbar_demux:src7_ready
	wire          cmd_xbar_demux_src8_endofpacket;                                                                                                  // cmd_xbar_demux:src8_endofpacket -> cmd_xbar_mux_008:sink0_endofpacket
	wire          cmd_xbar_demux_src8_valid;                                                                                                        // cmd_xbar_demux:src8_valid -> cmd_xbar_mux_008:sink0_valid
	wire          cmd_xbar_demux_src8_startofpacket;                                                                                                // cmd_xbar_demux:src8_startofpacket -> cmd_xbar_mux_008:sink0_startofpacket
	wire  [108:0] cmd_xbar_demux_src8_data;                                                                                                         // cmd_xbar_demux:src8_data -> cmd_xbar_mux_008:sink0_data
	wire   [18:0] cmd_xbar_demux_src8_channel;                                                                                                      // cmd_xbar_demux:src8_channel -> cmd_xbar_mux_008:sink0_channel
	wire          cmd_xbar_demux_src8_ready;                                                                                                        // cmd_xbar_mux_008:sink0_ready -> cmd_xbar_demux:src8_ready
	wire          cmd_xbar_demux_src9_endofpacket;                                                                                                  // cmd_xbar_demux:src9_endofpacket -> cmd_xbar_mux_009:sink0_endofpacket
	wire          cmd_xbar_demux_src9_valid;                                                                                                        // cmd_xbar_demux:src9_valid -> cmd_xbar_mux_009:sink0_valid
	wire          cmd_xbar_demux_src9_startofpacket;                                                                                                // cmd_xbar_demux:src9_startofpacket -> cmd_xbar_mux_009:sink0_startofpacket
	wire  [108:0] cmd_xbar_demux_src9_data;                                                                                                         // cmd_xbar_demux:src9_data -> cmd_xbar_mux_009:sink0_data
	wire   [18:0] cmd_xbar_demux_src9_channel;                                                                                                      // cmd_xbar_demux:src9_channel -> cmd_xbar_mux_009:sink0_channel
	wire          cmd_xbar_demux_src9_ready;                                                                                                        // cmd_xbar_mux_009:sink0_ready -> cmd_xbar_demux:src9_ready
	wire          cmd_xbar_demux_src10_endofpacket;                                                                                                 // cmd_xbar_demux:src10_endofpacket -> cmd_xbar_mux_010:sink0_endofpacket
	wire          cmd_xbar_demux_src10_valid;                                                                                                       // cmd_xbar_demux:src10_valid -> cmd_xbar_mux_010:sink0_valid
	wire          cmd_xbar_demux_src10_startofpacket;                                                                                               // cmd_xbar_demux:src10_startofpacket -> cmd_xbar_mux_010:sink0_startofpacket
	wire  [108:0] cmd_xbar_demux_src10_data;                                                                                                        // cmd_xbar_demux:src10_data -> cmd_xbar_mux_010:sink0_data
	wire   [18:0] cmd_xbar_demux_src10_channel;                                                                                                     // cmd_xbar_demux:src10_channel -> cmd_xbar_mux_010:sink0_channel
	wire          cmd_xbar_demux_src10_ready;                                                                                                       // cmd_xbar_mux_010:sink0_ready -> cmd_xbar_demux:src10_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                                              // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                                                    // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                                                            // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src0_data;                                                                                                     // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src0_channel;                                                                                                  // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                                                    // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                                              // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                                                    // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                                                            // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src1_data;                                                                                                     // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src1_channel;                                                                                                  // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                                                    // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                                                              // cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                                                    // cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                                                            // cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src3_data;                                                                                                     // cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src3_channel;                                                                                                  // cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	wire          cmd_xbar_demux_001_src3_ready;                                                                                                    // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                                                              // cmd_xbar_demux_001:src4_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                                                    // cmd_xbar_demux_001:src4_valid -> cmd_xbar_mux_004:sink1_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                                                            // cmd_xbar_demux_001:src4_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src4_data;                                                                                                     // cmd_xbar_demux_001:src4_data -> cmd_xbar_mux_004:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src4_channel;                                                                                                  // cmd_xbar_demux_001:src4_channel -> cmd_xbar_mux_004:sink1_channel
	wire          cmd_xbar_demux_001_src4_ready;                                                                                                    // cmd_xbar_mux_004:sink1_ready -> cmd_xbar_demux_001:src4_ready
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                                                              // cmd_xbar_demux_001:src5_endofpacket -> cmd_xbar_mux_005:sink1_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                                                    // cmd_xbar_demux_001:src5_valid -> cmd_xbar_mux_005:sink1_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                                                            // cmd_xbar_demux_001:src5_startofpacket -> cmd_xbar_mux_005:sink1_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src5_data;                                                                                                     // cmd_xbar_demux_001:src5_data -> cmd_xbar_mux_005:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src5_channel;                                                                                                  // cmd_xbar_demux_001:src5_channel -> cmd_xbar_mux_005:sink1_channel
	wire          cmd_xbar_demux_001_src5_ready;                                                                                                    // cmd_xbar_mux_005:sink1_ready -> cmd_xbar_demux_001:src5_ready
	wire          cmd_xbar_demux_001_src6_endofpacket;                                                                                              // cmd_xbar_demux_001:src6_endofpacket -> cmd_xbar_mux_006:sink1_endofpacket
	wire          cmd_xbar_demux_001_src6_valid;                                                                                                    // cmd_xbar_demux_001:src6_valid -> cmd_xbar_mux_006:sink1_valid
	wire          cmd_xbar_demux_001_src6_startofpacket;                                                                                            // cmd_xbar_demux_001:src6_startofpacket -> cmd_xbar_mux_006:sink1_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src6_data;                                                                                                     // cmd_xbar_demux_001:src6_data -> cmd_xbar_mux_006:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src6_channel;                                                                                                  // cmd_xbar_demux_001:src6_channel -> cmd_xbar_mux_006:sink1_channel
	wire          cmd_xbar_demux_001_src6_ready;                                                                                                    // cmd_xbar_mux_006:sink1_ready -> cmd_xbar_demux_001:src6_ready
	wire          cmd_xbar_demux_001_src7_endofpacket;                                                                                              // cmd_xbar_demux_001:src7_endofpacket -> cmd_xbar_mux_007:sink1_endofpacket
	wire          cmd_xbar_demux_001_src7_valid;                                                                                                    // cmd_xbar_demux_001:src7_valid -> cmd_xbar_mux_007:sink1_valid
	wire          cmd_xbar_demux_001_src7_startofpacket;                                                                                            // cmd_xbar_demux_001:src7_startofpacket -> cmd_xbar_mux_007:sink1_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src7_data;                                                                                                     // cmd_xbar_demux_001:src7_data -> cmd_xbar_mux_007:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src7_channel;                                                                                                  // cmd_xbar_demux_001:src7_channel -> cmd_xbar_mux_007:sink1_channel
	wire          cmd_xbar_demux_001_src7_ready;                                                                                                    // cmd_xbar_mux_007:sink1_ready -> cmd_xbar_demux_001:src7_ready
	wire          cmd_xbar_demux_001_src8_endofpacket;                                                                                              // cmd_xbar_demux_001:src8_endofpacket -> cmd_xbar_mux_008:sink1_endofpacket
	wire          cmd_xbar_demux_001_src8_valid;                                                                                                    // cmd_xbar_demux_001:src8_valid -> cmd_xbar_mux_008:sink1_valid
	wire          cmd_xbar_demux_001_src8_startofpacket;                                                                                            // cmd_xbar_demux_001:src8_startofpacket -> cmd_xbar_mux_008:sink1_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src8_data;                                                                                                     // cmd_xbar_demux_001:src8_data -> cmd_xbar_mux_008:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src8_channel;                                                                                                  // cmd_xbar_demux_001:src8_channel -> cmd_xbar_mux_008:sink1_channel
	wire          cmd_xbar_demux_001_src8_ready;                                                                                                    // cmd_xbar_mux_008:sink1_ready -> cmd_xbar_demux_001:src8_ready
	wire          cmd_xbar_demux_001_src9_endofpacket;                                                                                              // cmd_xbar_demux_001:src9_endofpacket -> cmd_xbar_mux_009:sink1_endofpacket
	wire          cmd_xbar_demux_001_src9_valid;                                                                                                    // cmd_xbar_demux_001:src9_valid -> cmd_xbar_mux_009:sink1_valid
	wire          cmd_xbar_demux_001_src9_startofpacket;                                                                                            // cmd_xbar_demux_001:src9_startofpacket -> cmd_xbar_mux_009:sink1_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src9_data;                                                                                                     // cmd_xbar_demux_001:src9_data -> cmd_xbar_mux_009:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src9_channel;                                                                                                  // cmd_xbar_demux_001:src9_channel -> cmd_xbar_mux_009:sink1_channel
	wire          cmd_xbar_demux_001_src9_ready;                                                                                                    // cmd_xbar_mux_009:sink1_ready -> cmd_xbar_demux_001:src9_ready
	wire          cmd_xbar_demux_001_src10_endofpacket;                                                                                             // cmd_xbar_demux_001:src10_endofpacket -> cmd_xbar_mux_010:sink1_endofpacket
	wire          cmd_xbar_demux_001_src10_valid;                                                                                                   // cmd_xbar_demux_001:src10_valid -> cmd_xbar_mux_010:sink1_valid
	wire          cmd_xbar_demux_001_src10_startofpacket;                                                                                           // cmd_xbar_demux_001:src10_startofpacket -> cmd_xbar_mux_010:sink1_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src10_data;                                                                                                    // cmd_xbar_demux_001:src10_data -> cmd_xbar_mux_010:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src10_channel;                                                                                                 // cmd_xbar_demux_001:src10_channel -> cmd_xbar_mux_010:sink1_channel
	wire          cmd_xbar_demux_001_src10_ready;                                                                                                   // cmd_xbar_mux_010:sink1_ready -> cmd_xbar_demux_001:src10_ready
	wire          cmd_xbar_demux_001_src12_endofpacket;                                                                                             // cmd_xbar_demux_001:src12_endofpacket -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src12_valid;                                                                                                   // cmd_xbar_demux_001:src12_valid -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src12_startofpacket;                                                                                           // cmd_xbar_demux_001:src12_startofpacket -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src12_data;                                                                                                    // cmd_xbar_demux_001:src12_data -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_demux_001_src12_channel;                                                                                                 // cmd_xbar_demux_001:src12_channel -> JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src13_endofpacket;                                                                                             // cmd_xbar_demux_001:src13_endofpacket -> video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src13_valid;                                                                                                   // cmd_xbar_demux_001:src13_valid -> video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src13_startofpacket;                                                                                           // cmd_xbar_demux_001:src13_startofpacket -> video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src13_data;                                                                                                    // cmd_xbar_demux_001:src13_data -> video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_demux_001_src13_channel;                                                                                                 // cmd_xbar_demux_001:src13_channel -> video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src14_endofpacket;                                                                                             // cmd_xbar_demux_001:src14_endofpacket -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src14_valid;                                                                                                   // cmd_xbar_demux_001:src14_valid -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src14_startofpacket;                                                                                           // cmd_xbar_demux_001:src14_startofpacket -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src14_data;                                                                                                    // cmd_xbar_demux_001:src14_data -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_demux_001_src14_channel;                                                                                                 // cmd_xbar_demux_001:src14_channel -> video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src17_endofpacket;                                                                                             // cmd_xbar_demux_001:src17_endofpacket -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src17_valid;                                                                                                   // cmd_xbar_demux_001:src17_valid -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src17_startofpacket;                                                                                           // cmd_xbar_demux_001:src17_startofpacket -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src17_data;                                                                                                    // cmd_xbar_demux_001:src17_data -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_demux_001_src17_channel;                                                                                                 // cmd_xbar_demux_001:src17_channel -> audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src18_endofpacket;                                                                                             // cmd_xbar_demux_001:src18_endofpacket -> cmd_xbar_mux_018:sink0_endofpacket
	wire          cmd_xbar_demux_001_src18_valid;                                                                                                   // cmd_xbar_demux_001:src18_valid -> cmd_xbar_mux_018:sink0_valid
	wire          cmd_xbar_demux_001_src18_startofpacket;                                                                                           // cmd_xbar_demux_001:src18_startofpacket -> cmd_xbar_mux_018:sink0_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src18_data;                                                                                                    // cmd_xbar_demux_001:src18_data -> cmd_xbar_mux_018:sink0_data
	wire   [18:0] cmd_xbar_demux_001_src18_channel;                                                                                                 // cmd_xbar_demux_001:src18_channel -> cmd_xbar_mux_018:sink0_channel
	wire          cmd_xbar_demux_001_src18_ready;                                                                                                   // cmd_xbar_mux_018:sink0_ready -> cmd_xbar_demux_001:src18_ready
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                                                              // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_016:sink1_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                                                    // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_016:sink1_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                                                            // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_016:sink1_startofpacket
	wire   [90:0] cmd_xbar_demux_002_src0_data;                                                                                                     // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_016:sink1_data
	wire   [18:0] cmd_xbar_demux_002_src0_channel;                                                                                                  // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_016:sink1_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                                                    // cmd_xbar_mux_016:sink1_ready -> cmd_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_src0_endofpacket;                                                                                                  // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                                                        // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                                                // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [108:0] rsp_xbar_demux_src0_data;                                                                                                         // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [18:0] rsp_xbar_demux_src0_channel;                                                                                                      // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                                                        // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                                                  // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                                                        // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                                                // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [108:0] rsp_xbar_demux_src1_data;                                                                                                         // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [18:0] rsp_xbar_demux_src1_channel;                                                                                                      // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                                                        // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                                              // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                                                    // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                                                            // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [108:0] rsp_xbar_demux_001_src0_data;                                                                                                     // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [18:0] rsp_xbar_demux_001_src0_channel;                                                                                                  // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                                                    // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                                                              // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                                                    // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                                                            // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [108:0] rsp_xbar_demux_001_src1_data;                                                                                                     // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [18:0] rsp_xbar_demux_001_src1_channel;                                                                                                  // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                                                    // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                                              // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                                                    // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                                                            // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [108:0] rsp_xbar_demux_003_src0_data;                                                                                                     // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire   [18:0] rsp_xbar_demux_003_src0_channel;                                                                                                  // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                                                    // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_003_src1_endofpacket;                                                                                              // rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_003_src1_valid;                                                                                                    // rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_003_src1_startofpacket;                                                                                            // rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [108:0] rsp_xbar_demux_003_src1_data;                                                                                                     // rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	wire   [18:0] rsp_xbar_demux_003_src1_channel;                                                                                                  // rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_003_src1_ready;                                                                                                    // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                                              // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                                                    // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                                                            // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire  [108:0] rsp_xbar_demux_004_src0_data;                                                                                                     // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	wire   [18:0] rsp_xbar_demux_004_src0_channel;                                                                                                  // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                                                    // rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_004_src1_endofpacket;                                                                                              // rsp_xbar_demux_004:src1_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_004_src1_valid;                                                                                                    // rsp_xbar_demux_004:src1_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_004_src1_startofpacket;                                                                                            // rsp_xbar_demux_004:src1_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [108:0] rsp_xbar_demux_004_src1_data;                                                                                                     // rsp_xbar_demux_004:src1_data -> rsp_xbar_mux_001:sink4_data
	wire   [18:0] rsp_xbar_demux_004_src1_channel;                                                                                                  // rsp_xbar_demux_004:src1_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_004_src1_ready;                                                                                                    // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src1_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                                              // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux:sink5_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                                                    // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux:sink5_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                                                            // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux:sink5_startofpacket
	wire  [108:0] rsp_xbar_demux_005_src0_data;                                                                                                     // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux:sink5_data
	wire   [18:0] rsp_xbar_demux_005_src0_channel;                                                                                                  // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux:sink5_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                                                    // rsp_xbar_mux:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_005_src1_endofpacket;                                                                                              // rsp_xbar_demux_005:src1_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          rsp_xbar_demux_005_src1_valid;                                                                                                    // rsp_xbar_demux_005:src1_valid -> rsp_xbar_mux_001:sink5_valid
	wire          rsp_xbar_demux_005_src1_startofpacket;                                                                                            // rsp_xbar_demux_005:src1_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [108:0] rsp_xbar_demux_005_src1_data;                                                                                                     // rsp_xbar_demux_005:src1_data -> rsp_xbar_mux_001:sink5_data
	wire   [18:0] rsp_xbar_demux_005_src1_channel;                                                                                                  // rsp_xbar_demux_005:src1_channel -> rsp_xbar_mux_001:sink5_channel
	wire          rsp_xbar_demux_005_src1_ready;                                                                                                    // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src1_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                                              // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux:sink6_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                                                    // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux:sink6_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                                                            // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux:sink6_startofpacket
	wire  [108:0] rsp_xbar_demux_006_src0_data;                                                                                                     // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux:sink6_data
	wire   [18:0] rsp_xbar_demux_006_src0_channel;                                                                                                  // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux:sink6_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                                                    // rsp_xbar_mux:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_006_src1_endofpacket;                                                                                              // rsp_xbar_demux_006:src1_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire          rsp_xbar_demux_006_src1_valid;                                                                                                    // rsp_xbar_demux_006:src1_valid -> rsp_xbar_mux_001:sink6_valid
	wire          rsp_xbar_demux_006_src1_startofpacket;                                                                                            // rsp_xbar_demux_006:src1_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [108:0] rsp_xbar_demux_006_src1_data;                                                                                                     // rsp_xbar_demux_006:src1_data -> rsp_xbar_mux_001:sink6_data
	wire   [18:0] rsp_xbar_demux_006_src1_channel;                                                                                                  // rsp_xbar_demux_006:src1_channel -> rsp_xbar_mux_001:sink6_channel
	wire          rsp_xbar_demux_006_src1_ready;                                                                                                    // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src1_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                                              // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux:sink7_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                                                    // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux:sink7_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                                                            // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux:sink7_startofpacket
	wire  [108:0] rsp_xbar_demux_007_src0_data;                                                                                                     // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux:sink7_data
	wire   [18:0] rsp_xbar_demux_007_src0_channel;                                                                                                  // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux:sink7_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                                                    // rsp_xbar_mux:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_007_src1_endofpacket;                                                                                              // rsp_xbar_demux_007:src1_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire          rsp_xbar_demux_007_src1_valid;                                                                                                    // rsp_xbar_demux_007:src1_valid -> rsp_xbar_mux_001:sink7_valid
	wire          rsp_xbar_demux_007_src1_startofpacket;                                                                                            // rsp_xbar_demux_007:src1_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [108:0] rsp_xbar_demux_007_src1_data;                                                                                                     // rsp_xbar_demux_007:src1_data -> rsp_xbar_mux_001:sink7_data
	wire   [18:0] rsp_xbar_demux_007_src1_channel;                                                                                                  // rsp_xbar_demux_007:src1_channel -> rsp_xbar_mux_001:sink7_channel
	wire          rsp_xbar_demux_007_src1_ready;                                                                                                    // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src1_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                                              // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux:sink8_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                                                    // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux:sink8_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                                                            // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux:sink8_startofpacket
	wire  [108:0] rsp_xbar_demux_008_src0_data;                                                                                                     // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux:sink8_data
	wire   [18:0] rsp_xbar_demux_008_src0_channel;                                                                                                  // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux:sink8_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                                                    // rsp_xbar_mux:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire          rsp_xbar_demux_008_src1_endofpacket;                                                                                              // rsp_xbar_demux_008:src1_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire          rsp_xbar_demux_008_src1_valid;                                                                                                    // rsp_xbar_demux_008:src1_valid -> rsp_xbar_mux_001:sink8_valid
	wire          rsp_xbar_demux_008_src1_startofpacket;                                                                                            // rsp_xbar_demux_008:src1_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [108:0] rsp_xbar_demux_008_src1_data;                                                                                                     // rsp_xbar_demux_008:src1_data -> rsp_xbar_mux_001:sink8_data
	wire   [18:0] rsp_xbar_demux_008_src1_channel;                                                                                                  // rsp_xbar_demux_008:src1_channel -> rsp_xbar_mux_001:sink8_channel
	wire          rsp_xbar_demux_008_src1_ready;                                                                                                    // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src1_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                                              // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux:sink9_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                                                    // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux:sink9_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                                                            // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux:sink9_startofpacket
	wire  [108:0] rsp_xbar_demux_009_src0_data;                                                                                                     // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux:sink9_data
	wire   [18:0] rsp_xbar_demux_009_src0_channel;                                                                                                  // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux:sink9_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                                                    // rsp_xbar_mux:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_009_src1_endofpacket;                                                                                              // rsp_xbar_demux_009:src1_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire          rsp_xbar_demux_009_src1_valid;                                                                                                    // rsp_xbar_demux_009:src1_valid -> rsp_xbar_mux_001:sink9_valid
	wire          rsp_xbar_demux_009_src1_startofpacket;                                                                                            // rsp_xbar_demux_009:src1_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [108:0] rsp_xbar_demux_009_src1_data;                                                                                                     // rsp_xbar_demux_009:src1_data -> rsp_xbar_mux_001:sink9_data
	wire   [18:0] rsp_xbar_demux_009_src1_channel;                                                                                                  // rsp_xbar_demux_009:src1_channel -> rsp_xbar_mux_001:sink9_channel
	wire          rsp_xbar_demux_009_src1_ready;                                                                                                    // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src1_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                                              // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux:sink10_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                                                    // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux:sink10_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                                                            // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux:sink10_startofpacket
	wire  [108:0] rsp_xbar_demux_010_src0_data;                                                                                                     // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux:sink10_data
	wire   [18:0] rsp_xbar_demux_010_src0_channel;                                                                                                  // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux:sink10_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                                                    // rsp_xbar_mux:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire          rsp_xbar_demux_010_src1_endofpacket;                                                                                              // rsp_xbar_demux_010:src1_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire          rsp_xbar_demux_010_src1_valid;                                                                                                    // rsp_xbar_demux_010:src1_valid -> rsp_xbar_mux_001:sink10_valid
	wire          rsp_xbar_demux_010_src1_startofpacket;                                                                                            // rsp_xbar_demux_010:src1_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [108:0] rsp_xbar_demux_010_src1_data;                                                                                                     // rsp_xbar_demux_010:src1_data -> rsp_xbar_mux_001:sink10_data
	wire   [18:0] rsp_xbar_demux_010_src1_channel;                                                                                                  // rsp_xbar_demux_010:src1_channel -> rsp_xbar_mux_001:sink10_channel
	wire          rsp_xbar_demux_010_src1_ready;                                                                                                    // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src1_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                                                              // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                                                    // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_001:sink12_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                                                            // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	wire  [108:0] rsp_xbar_demux_012_src0_data;                                                                                                     // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_001:sink12_data
	wire   [18:0] rsp_xbar_demux_012_src0_channel;                                                                                                  // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_001:sink12_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                                                    // rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                                                              // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                                                    // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_001:sink13_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                                                            // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	wire  [108:0] rsp_xbar_demux_013_src0_data;                                                                                                     // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_001:sink13_data
	wire   [18:0] rsp_xbar_demux_013_src0_channel;                                                                                                  // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_001:sink13_channel
	wire          rsp_xbar_demux_013_src0_ready;                                                                                                    // rsp_xbar_mux_001:sink13_ready -> rsp_xbar_demux_013:src0_ready
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                                                              // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_001:sink14_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                                                    // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_001:sink14_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                                                            // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_001:sink14_startofpacket
	wire  [108:0] rsp_xbar_demux_014_src0_data;                                                                                                     // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_001:sink14_data
	wire   [18:0] rsp_xbar_demux_014_src0_channel;                                                                                                  // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_001:sink14_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                                                    // rsp_xbar_mux_001:sink14_ready -> rsp_xbar_demux_014:src0_ready
	wire          rsp_xbar_demux_016_src1_endofpacket;                                                                                              // rsp_xbar_demux_016:src1_endofpacket -> rsp_xbar_mux_002:sink0_endofpacket
	wire          rsp_xbar_demux_016_src1_valid;                                                                                                    // rsp_xbar_demux_016:src1_valid -> rsp_xbar_mux_002:sink0_valid
	wire          rsp_xbar_demux_016_src1_startofpacket;                                                                                            // rsp_xbar_demux_016:src1_startofpacket -> rsp_xbar_mux_002:sink0_startofpacket
	wire   [90:0] rsp_xbar_demux_016_src1_data;                                                                                                     // rsp_xbar_demux_016:src1_data -> rsp_xbar_mux_002:sink0_data
	wire   [18:0] rsp_xbar_demux_016_src1_channel;                                                                                                  // rsp_xbar_demux_016:src1_channel -> rsp_xbar_mux_002:sink0_channel
	wire          rsp_xbar_demux_016_src1_ready;                                                                                                    // rsp_xbar_mux_002:sink0_ready -> rsp_xbar_demux_016:src1_ready
	wire          rsp_xbar_demux_017_src0_endofpacket;                                                                                              // rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux_001:sink17_endofpacket
	wire          rsp_xbar_demux_017_src0_valid;                                                                                                    // rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux_001:sink17_valid
	wire          rsp_xbar_demux_017_src0_startofpacket;                                                                                            // rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux_001:sink17_startofpacket
	wire  [108:0] rsp_xbar_demux_017_src0_data;                                                                                                     // rsp_xbar_demux_017:src0_data -> rsp_xbar_mux_001:sink17_data
	wire   [18:0] rsp_xbar_demux_017_src0_channel;                                                                                                  // rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux_001:sink17_channel
	wire          rsp_xbar_demux_017_src0_ready;                                                                                                    // rsp_xbar_mux_001:sink17_ready -> rsp_xbar_demux_017:src0_ready
	wire          rsp_xbar_demux_018_src0_endofpacket;                                                                                              // rsp_xbar_demux_018:src0_endofpacket -> rsp_xbar_mux_001:sink18_endofpacket
	wire          rsp_xbar_demux_018_src0_valid;                                                                                                    // rsp_xbar_demux_018:src0_valid -> rsp_xbar_mux_001:sink18_valid
	wire          rsp_xbar_demux_018_src0_startofpacket;                                                                                            // rsp_xbar_demux_018:src0_startofpacket -> rsp_xbar_mux_001:sink18_startofpacket
	wire  [108:0] rsp_xbar_demux_018_src0_data;                                                                                                     // rsp_xbar_demux_018:src0_data -> rsp_xbar_mux_001:sink18_data
	wire   [18:0] rsp_xbar_demux_018_src0_channel;                                                                                                  // rsp_xbar_demux_018:src0_channel -> rsp_xbar_mux_001:sink18_channel
	wire          rsp_xbar_demux_018_src0_ready;                                                                                                    // rsp_xbar_mux_001:sink18_ready -> rsp_xbar_demux_018:src0_ready
	wire          limiter_cmd_src_endofpacket;                                                                                                      // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                                                    // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [108:0] limiter_cmd_src_data;                                                                                                             // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire   [18:0] limiter_cmd_src_channel;                                                                                                          // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_cmd_src_ready;                                                                                                            // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                                                     // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                                                           // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                                                   // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [108:0] rsp_xbar_mux_src_data;                                                                                                            // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire   [18:0] rsp_xbar_mux_src_channel;                                                                                                         // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_src_ready;                                                                                                           // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire          limiter_001_cmd_src_endofpacket;                                                                                                  // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          limiter_001_cmd_src_startofpacket;                                                                                                // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [108:0] limiter_001_cmd_src_data;                                                                                                         // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire   [18:0] limiter_001_cmd_src_channel;                                                                                                      // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire          limiter_001_cmd_src_ready;                                                                                                        // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                                                 // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                                                       // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                                               // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [108:0] rsp_xbar_mux_001_src_data;                                                                                                        // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire   [18:0] rsp_xbar_mux_001_src_channel;                                                                                                     // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                                                       // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire          limiter_002_cmd_src_endofpacket;                                                                                                  // limiter_002:cmd_src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          limiter_002_cmd_src_startofpacket;                                                                                                // limiter_002:cmd_src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire   [90:0] limiter_002_cmd_src_data;                                                                                                         // limiter_002:cmd_src_data -> cmd_xbar_demux_002:sink_data
	wire   [18:0] limiter_002_cmd_src_channel;                                                                                                      // limiter_002:cmd_src_channel -> cmd_xbar_demux_002:sink_channel
	wire          limiter_002_cmd_src_ready;                                                                                                        // cmd_xbar_demux_002:sink_ready -> limiter_002:cmd_src_ready
	wire          rsp_xbar_mux_002_src_endofpacket;                                                                                                 // rsp_xbar_mux_002:src_endofpacket -> limiter_002:rsp_sink_endofpacket
	wire          rsp_xbar_mux_002_src_valid;                                                                                                       // rsp_xbar_mux_002:src_valid -> limiter_002:rsp_sink_valid
	wire          rsp_xbar_mux_002_src_startofpacket;                                                                                               // rsp_xbar_mux_002:src_startofpacket -> limiter_002:rsp_sink_startofpacket
	wire   [90:0] rsp_xbar_mux_002_src_data;                                                                                                        // rsp_xbar_mux_002:src_data -> limiter_002:rsp_sink_data
	wire   [18:0] rsp_xbar_mux_002_src_channel;                                                                                                     // rsp_xbar_mux_002:src_channel -> limiter_002:rsp_sink_channel
	wire          rsp_xbar_mux_002_src_ready;                                                                                                       // limiter_002:rsp_sink_ready -> rsp_xbar_mux_002:src_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                                                     // cmd_xbar_mux:src_endofpacket -> nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                                                           // cmd_xbar_mux:src_valid -> nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                                                   // cmd_xbar_mux:src_startofpacket -> nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_mux_src_data;                                                                                                            // cmd_xbar_mux:src_data -> nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_src_channel;                                                                                                         // cmd_xbar_mux:src_channel -> nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                                                           // nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                                                        // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                                              // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                                                      // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [108:0] id_router_src_data;                                                                                                               // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [18:0] id_router_src_channel;                                                                                                            // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                                              // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                                                 // cmd_xbar_mux_001:src_endofpacket -> onchip_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                                                       // cmd_xbar_mux_001:src_valid -> onchip_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                                               // cmd_xbar_mux_001:src_startofpacket -> onchip_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_mux_001_src_data;                                                                                                        // cmd_xbar_mux_001:src_data -> onchip_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_001_src_channel;                                                                                                     // cmd_xbar_mux_001:src_channel -> onchip_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                                                       // onchip_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire          id_router_001_src_endofpacket;                                                                                                    // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                                                          // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                                                  // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [108:0] id_router_001_src_data;                                                                                                           // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [18:0] id_router_001_src_channel;                                                                                                        // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                                                          // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_mux_002_src_endofpacket;                                                                                                 // cmd_xbar_mux_002:src_endofpacket -> burst_adapter:sink0_endofpacket
	wire          cmd_xbar_mux_002_src_valid;                                                                                                       // cmd_xbar_mux_002:src_valid -> burst_adapter:sink0_valid
	wire          cmd_xbar_mux_002_src_startofpacket;                                                                                               // cmd_xbar_mux_002:src_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [90:0] cmd_xbar_mux_002_src_data;                                                                                                        // cmd_xbar_mux_002:src_data -> burst_adapter:sink0_data
	wire   [18:0] cmd_xbar_mux_002_src_channel;                                                                                                     // cmd_xbar_mux_002:src_channel -> burst_adapter:sink0_channel
	wire          cmd_xbar_mux_002_src_ready;                                                                                                       // burst_adapter:sink0_ready -> cmd_xbar_mux_002:src_ready
	wire          id_router_002_src_endofpacket;                                                                                                    // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                                                          // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                                                  // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire   [90:0] id_router_002_src_data;                                                                                                           // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [18:0] id_router_002_src_channel;                                                                                                        // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                                                          // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_mux_003_src_endofpacket;                                                                                                 // cmd_xbar_mux_003:src_endofpacket -> LEDG_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_003_src_valid;                                                                                                       // cmd_xbar_mux_003:src_valid -> LEDG_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_003_src_startofpacket;                                                                                               // cmd_xbar_mux_003:src_startofpacket -> LEDG_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_mux_003_src_data;                                                                                                        // cmd_xbar_mux_003:src_data -> LEDG_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_003_src_channel;                                                                                                     // cmd_xbar_mux_003:src_channel -> LEDG_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_003_src_ready;                                                                                                       // LEDG_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_003:src_ready
	wire          id_router_003_src_endofpacket;                                                                                                    // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                                                          // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                                                  // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [108:0] id_router_003_src_data;                                                                                                           // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [18:0] id_router_003_src_channel;                                                                                                        // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                                                          // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_mux_004_src_endofpacket;                                                                                                 // cmd_xbar_mux_004:src_endofpacket -> LEDR_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_004_src_valid;                                                                                                       // cmd_xbar_mux_004:src_valid -> LEDR_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_004_src_startofpacket;                                                                                               // cmd_xbar_mux_004:src_startofpacket -> LEDR_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_mux_004_src_data;                                                                                                        // cmd_xbar_mux_004:src_data -> LEDR_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_004_src_channel;                                                                                                     // cmd_xbar_mux_004:src_channel -> LEDR_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_004_src_ready;                                                                                                       // LEDR_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_004:src_ready
	wire          id_router_004_src_endofpacket;                                                                                                    // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                                                          // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                                                  // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [108:0] id_router_004_src_data;                                                                                                           // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [18:0] id_router_004_src_channel;                                                                                                        // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                                                          // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_mux_005_src_endofpacket;                                                                                                 // cmd_xbar_mux_005:src_endofpacket -> switches_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_005_src_valid;                                                                                                       // cmd_xbar_mux_005:src_valid -> switches_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_005_src_startofpacket;                                                                                               // cmd_xbar_mux_005:src_startofpacket -> switches_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_mux_005_src_data;                                                                                                        // cmd_xbar_mux_005:src_data -> switches_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_005_src_channel;                                                                                                     // cmd_xbar_mux_005:src_channel -> switches_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_005_src_ready;                                                                                                       // switches_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_005:src_ready
	wire          id_router_005_src_endofpacket;                                                                                                    // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                                                          // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                                                  // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [108:0] id_router_005_src_data;                                                                                                           // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [18:0] id_router_005_src_channel;                                                                                                        // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                                                          // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_mux_006_src_endofpacket;                                                                                                 // cmd_xbar_mux_006:src_endofpacket -> key_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_006_src_valid;                                                                                                       // cmd_xbar_mux_006:src_valid -> key_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_006_src_startofpacket;                                                                                               // cmd_xbar_mux_006:src_startofpacket -> key_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_mux_006_src_data;                                                                                                        // cmd_xbar_mux_006:src_data -> key_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_006_src_channel;                                                                                                     // cmd_xbar_mux_006:src_channel -> key_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_006_src_ready;                                                                                                       // key_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_006:src_ready
	wire          id_router_006_src_endofpacket;                                                                                                    // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                                                          // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                                                  // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [108:0] id_router_006_src_data;                                                                                                           // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [18:0] id_router_006_src_channel;                                                                                                        // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                                                          // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_mux_007_src_endofpacket;                                                                                                 // cmd_xbar_mux_007:src_endofpacket -> sdcard_timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_007_src_valid;                                                                                                       // cmd_xbar_mux_007:src_valid -> sdcard_timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_007_src_startofpacket;                                                                                               // cmd_xbar_mux_007:src_startofpacket -> sdcard_timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_mux_007_src_data;                                                                                                        // cmd_xbar_mux_007:src_data -> sdcard_timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_007_src_channel;                                                                                                     // cmd_xbar_mux_007:src_channel -> sdcard_timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_007_src_ready;                                                                                                       // sdcard_timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_007:src_ready
	wire          id_router_007_src_endofpacket;                                                                                                    // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                                                          // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                                                  // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [108:0] id_router_007_src_data;                                                                                                           // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [18:0] id_router_007_src_channel;                                                                                                        // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                                                          // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_mux_008_src_endofpacket;                                                                                                 // cmd_xbar_mux_008:src_endofpacket -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_008_src_valid;                                                                                                       // cmd_xbar_mux_008:src_valid -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_008_src_startofpacket;                                                                                               // cmd_xbar_mux_008:src_startofpacket -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_mux_008_src_data;                                                                                                        // cmd_xbar_mux_008:src_data -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_008_src_channel;                                                                                                     // cmd_xbar_mux_008:src_channel -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_008_src_ready;                                                                                                       // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_008:src_ready
	wire          id_router_008_src_endofpacket;                                                                                                    // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                                                          // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                                                  // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [108:0] id_router_008_src_data;                                                                                                           // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [18:0] id_router_008_src_channel;                                                                                                        // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                                                          // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_mux_009_src_endofpacket;                                                                                                 // cmd_xbar_mux_009:src_endofpacket -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_009_src_valid;                                                                                                       // cmd_xbar_mux_009:src_valid -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_009_src_startofpacket;                                                                                               // cmd_xbar_mux_009:src_startofpacket -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_mux_009_src_data;                                                                                                        // cmd_xbar_mux_009:src_data -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_009_src_channel;                                                                                                     // cmd_xbar_mux_009:src_channel -> ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_009_src_ready;                                                                                                       // ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_009:src_ready
	wire          id_router_009_src_endofpacket;                                                                                                    // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                                                          // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                                                  // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [108:0] id_router_009_src_data;                                                                                                           // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [18:0] id_router_009_src_channel;                                                                                                        // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                                                          // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_mux_010_src_endofpacket;                                                                                                 // cmd_xbar_mux_010:src_endofpacket -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_010_src_valid;                                                                                                       // cmd_xbar_mux_010:src_valid -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_010_src_startofpacket;                                                                                               // cmd_xbar_mux_010:src_startofpacket -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_mux_010_src_data;                                                                                                        // cmd_xbar_mux_010:src_data -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_010_src_channel;                                                                                                     // cmd_xbar_mux_010:src_channel -> audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_010_src_ready;                                                                                                       // audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_010:src_ready
	wire          id_router_010_src_endofpacket;                                                                                                    // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                                                          // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                                                  // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [108:0] id_router_010_src_data;                                                                                                           // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [18:0] id_router_010_src_channel;                                                                                                        // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                                                          // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          width_adapter_002_src_ready;                                                                                                      // burst_adapter_001:sink0_ready -> width_adapter_002:out_ready
	wire          id_router_011_src_endofpacket;                                                                                                    // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                                                          // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                                                  // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire   [81:0] id_router_011_src_data;                                                                                                           // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire   [18:0] id_router_011_src_channel;                                                                                                        // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                                                          // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          cmd_xbar_demux_001_src12_ready;                                                                                                   // JTAG_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src12_ready
	wire          id_router_012_src_endofpacket;                                                                                                    // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                                                          // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                                                  // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [108:0] id_router_012_src_data;                                                                                                           // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire   [18:0] id_router_012_src_channel;                                                                                                        // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                                                          // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          cmd_xbar_demux_001_src13_ready;                                                                                                   // video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src13_ready
	wire          id_router_013_src_endofpacket;                                                                                                    // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                                                          // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                                                  // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [108:0] id_router_013_src_data;                                                                                                           // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire   [18:0] id_router_013_src_channel;                                                                                                        // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                                                          // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          cmd_xbar_demux_001_src14_ready;                                                                                                   // video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src14_ready
	wire          id_router_014_src_endofpacket;                                                                                                    // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          id_router_014_src_valid;                                                                                                          // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire          id_router_014_src_startofpacket;                                                                                                  // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [108:0] id_router_014_src_data;                                                                                                           // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire   [18:0] id_router_014_src_channel;                                                                                                        // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire          id_router_014_src_ready;                                                                                                          // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire          width_adapter_003_src_ready;                                                                                                      // burst_adapter_002:sink0_ready -> width_adapter_003:out_ready
	wire          id_router_015_src_endofpacket;                                                                                                    // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                                                          // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                                                  // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire   [81:0] id_router_015_src_data;                                                                                                           // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire   [18:0] id_router_015_src_channel;                                                                                                        // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                                                          // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire          cmd_xbar_mux_016_src_endofpacket;                                                                                                 // cmd_xbar_mux_016:src_endofpacket -> burst_adapter_003:sink0_endofpacket
	wire          cmd_xbar_mux_016_src_valid;                                                                                                       // cmd_xbar_mux_016:src_valid -> burst_adapter_003:sink0_valid
	wire          cmd_xbar_mux_016_src_startofpacket;                                                                                               // cmd_xbar_mux_016:src_startofpacket -> burst_adapter_003:sink0_startofpacket
	wire   [90:0] cmd_xbar_mux_016_src_data;                                                                                                        // cmd_xbar_mux_016:src_data -> burst_adapter_003:sink0_data
	wire   [18:0] cmd_xbar_mux_016_src_channel;                                                                                                     // cmd_xbar_mux_016:src_channel -> burst_adapter_003:sink0_channel
	wire          cmd_xbar_mux_016_src_ready;                                                                                                       // burst_adapter_003:sink0_ready -> cmd_xbar_mux_016:src_ready
	wire          id_router_016_src_endofpacket;                                                                                                    // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire          id_router_016_src_valid;                                                                                                          // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire          id_router_016_src_startofpacket;                                                                                                  // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire   [90:0] id_router_016_src_data;                                                                                                           // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire   [18:0] id_router_016_src_channel;                                                                                                        // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire          id_router_016_src_ready;                                                                                                          // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire          cmd_xbar_demux_001_src17_ready;                                                                                                   // audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src17_ready
	wire          id_router_017_src_endofpacket;                                                                                                    // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire          id_router_017_src_valid;                                                                                                          // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire          id_router_017_src_startofpacket;                                                                                                  // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire  [108:0] id_router_017_src_data;                                                                                                           // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire   [18:0] id_router_017_src_channel;                                                                                                        // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire          id_router_017_src_ready;                                                                                                          // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire          cmd_xbar_mux_018_src_endofpacket;                                                                                                 // cmd_xbar_mux_018:src_endofpacket -> usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_018_src_valid;                                                                                                       // cmd_xbar_mux_018:src_valid -> usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_018_src_startofpacket;                                                                                               // cmd_xbar_mux_018:src_startofpacket -> usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_mux_018_src_data;                                                                                                        // cmd_xbar_mux_018:src_data -> usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_018_src_channel;                                                                                                     // cmd_xbar_mux_018:src_channel -> usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_018_src_ready;                                                                                                       // usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_018:src_ready
	wire          id_router_018_src_endofpacket;                                                                                                    // id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire          id_router_018_src_valid;                                                                                                          // id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	wire          id_router_018_src_startofpacket;                                                                                                  // id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire  [108:0] id_router_018_src_data;                                                                                                           // id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	wire   [18:0] id_router_018_src_channel;                                                                                                        // id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	wire          id_router_018_src_ready;                                                                                                          // rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	wire          cmd_xbar_demux_src2_endofpacket;                                                                                                  // cmd_xbar_demux:src2_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                                                        // cmd_xbar_demux:src2_valid -> width_adapter:in_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                                                // cmd_xbar_demux:src2_startofpacket -> width_adapter:in_startofpacket
	wire  [108:0] cmd_xbar_demux_src2_data;                                                                                                         // cmd_xbar_demux:src2_data -> width_adapter:in_data
	wire   [18:0] cmd_xbar_demux_src2_channel;                                                                                                      // cmd_xbar_demux:src2_channel -> width_adapter:in_channel
	wire          cmd_xbar_demux_src2_ready;                                                                                                        // width_adapter:in_ready -> cmd_xbar_demux:src2_ready
	wire          width_adapter_src_endofpacket;                                                                                                    // width_adapter:out_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                                                          // width_adapter:out_valid -> cmd_xbar_mux_002:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                                                  // width_adapter:out_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire   [90:0] width_adapter_src_data;                                                                                                           // width_adapter:out_data -> cmd_xbar_mux_002:sink0_data
	wire          width_adapter_src_ready;                                                                                                          // cmd_xbar_mux_002:sink0_ready -> width_adapter:out_ready
	wire   [18:0] width_adapter_src_channel;                                                                                                        // width_adapter:out_channel -> cmd_xbar_mux_002:sink0_channel
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                                              // cmd_xbar_demux_001:src2_endofpacket -> width_adapter_001:in_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                                                    // cmd_xbar_demux_001:src2_valid -> width_adapter_001:in_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                                                            // cmd_xbar_demux_001:src2_startofpacket -> width_adapter_001:in_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src2_data;                                                                                                     // cmd_xbar_demux_001:src2_data -> width_adapter_001:in_data
	wire   [18:0] cmd_xbar_demux_001_src2_channel;                                                                                                  // cmd_xbar_demux_001:src2_channel -> width_adapter_001:in_channel
	wire          cmd_xbar_demux_001_src2_ready;                                                                                                    // width_adapter_001:in_ready -> cmd_xbar_demux_001:src2_ready
	wire          width_adapter_001_src_endofpacket;                                                                                                // width_adapter_001:out_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire          width_adapter_001_src_valid;                                                                                                      // width_adapter_001:out_valid -> cmd_xbar_mux_002:sink1_valid
	wire          width_adapter_001_src_startofpacket;                                                                                              // width_adapter_001:out_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire   [90:0] width_adapter_001_src_data;                                                                                                       // width_adapter_001:out_data -> cmd_xbar_mux_002:sink1_data
	wire          width_adapter_001_src_ready;                                                                                                      // cmd_xbar_mux_002:sink1_ready -> width_adapter_001:out_ready
	wire   [18:0] width_adapter_001_src_channel;                                                                                                    // width_adapter_001:out_channel -> cmd_xbar_mux_002:sink1_channel
	wire          cmd_xbar_demux_001_src11_endofpacket;                                                                                             // cmd_xbar_demux_001:src11_endofpacket -> width_adapter_002:in_endofpacket
	wire          cmd_xbar_demux_001_src11_valid;                                                                                                   // cmd_xbar_demux_001:src11_valid -> width_adapter_002:in_valid
	wire          cmd_xbar_demux_001_src11_startofpacket;                                                                                           // cmd_xbar_demux_001:src11_startofpacket -> width_adapter_002:in_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src11_data;                                                                                                    // cmd_xbar_demux_001:src11_data -> width_adapter_002:in_data
	wire   [18:0] cmd_xbar_demux_001_src11_channel;                                                                                                 // cmd_xbar_demux_001:src11_channel -> width_adapter_002:in_channel
	wire          cmd_xbar_demux_001_src11_ready;                                                                                                   // width_adapter_002:in_ready -> cmd_xbar_demux_001:src11_ready
	wire          width_adapter_002_src_endofpacket;                                                                                                // width_adapter_002:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire          width_adapter_002_src_valid;                                                                                                      // width_adapter_002:out_valid -> burst_adapter_001:sink0_valid
	wire          width_adapter_002_src_startofpacket;                                                                                              // width_adapter_002:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire   [81:0] width_adapter_002_src_data;                                                                                                       // width_adapter_002:out_data -> burst_adapter_001:sink0_data
	wire   [18:0] width_adapter_002_src_channel;                                                                                                    // width_adapter_002:out_channel -> burst_adapter_001:sink0_channel
	wire          cmd_xbar_demux_001_src15_endofpacket;                                                                                             // cmd_xbar_demux_001:src15_endofpacket -> width_adapter_003:in_endofpacket
	wire          cmd_xbar_demux_001_src15_valid;                                                                                                   // cmd_xbar_demux_001:src15_valid -> width_adapter_003:in_valid
	wire          cmd_xbar_demux_001_src15_startofpacket;                                                                                           // cmd_xbar_demux_001:src15_startofpacket -> width_adapter_003:in_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src15_data;                                                                                                    // cmd_xbar_demux_001:src15_data -> width_adapter_003:in_data
	wire   [18:0] cmd_xbar_demux_001_src15_channel;                                                                                                 // cmd_xbar_demux_001:src15_channel -> width_adapter_003:in_channel
	wire          cmd_xbar_demux_001_src15_ready;                                                                                                   // width_adapter_003:in_ready -> cmd_xbar_demux_001:src15_ready
	wire          width_adapter_003_src_endofpacket;                                                                                                // width_adapter_003:out_endofpacket -> burst_adapter_002:sink0_endofpacket
	wire          width_adapter_003_src_valid;                                                                                                      // width_adapter_003:out_valid -> burst_adapter_002:sink0_valid
	wire          width_adapter_003_src_startofpacket;                                                                                              // width_adapter_003:out_startofpacket -> burst_adapter_002:sink0_startofpacket
	wire   [81:0] width_adapter_003_src_data;                                                                                                       // width_adapter_003:out_data -> burst_adapter_002:sink0_data
	wire   [18:0] width_adapter_003_src_channel;                                                                                                    // width_adapter_003:out_channel -> burst_adapter_002:sink0_channel
	wire          cmd_xbar_demux_001_src16_endofpacket;                                                                                             // cmd_xbar_demux_001:src16_endofpacket -> width_adapter_004:in_endofpacket
	wire          cmd_xbar_demux_001_src16_valid;                                                                                                   // cmd_xbar_demux_001:src16_valid -> width_adapter_004:in_valid
	wire          cmd_xbar_demux_001_src16_startofpacket;                                                                                           // cmd_xbar_demux_001:src16_startofpacket -> width_adapter_004:in_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src16_data;                                                                                                    // cmd_xbar_demux_001:src16_data -> width_adapter_004:in_data
	wire   [18:0] cmd_xbar_demux_001_src16_channel;                                                                                                 // cmd_xbar_demux_001:src16_channel -> width_adapter_004:in_channel
	wire          cmd_xbar_demux_001_src16_ready;                                                                                                   // width_adapter_004:in_ready -> cmd_xbar_demux_001:src16_ready
	wire          width_adapter_004_src_endofpacket;                                                                                                // width_adapter_004:out_endofpacket -> cmd_xbar_mux_016:sink0_endofpacket
	wire          width_adapter_004_src_valid;                                                                                                      // width_adapter_004:out_valid -> cmd_xbar_mux_016:sink0_valid
	wire          width_adapter_004_src_startofpacket;                                                                                              // width_adapter_004:out_startofpacket -> cmd_xbar_mux_016:sink0_startofpacket
	wire   [90:0] width_adapter_004_src_data;                                                                                                       // width_adapter_004:out_data -> cmd_xbar_mux_016:sink0_data
	wire          width_adapter_004_src_ready;                                                                                                      // cmd_xbar_mux_016:sink0_ready -> width_adapter_004:out_ready
	wire   [18:0] width_adapter_004_src_channel;                                                                                                    // width_adapter_004:out_channel -> cmd_xbar_mux_016:sink0_channel
	wire          cmd_xbar_demux_002_src1_endofpacket;                                                                                              // cmd_xbar_demux_002:src1_endofpacket -> width_adapter_005:in_endofpacket
	wire          cmd_xbar_demux_002_src1_valid;                                                                                                    // cmd_xbar_demux_002:src1_valid -> width_adapter_005:in_valid
	wire          cmd_xbar_demux_002_src1_startofpacket;                                                                                            // cmd_xbar_demux_002:src1_startofpacket -> width_adapter_005:in_startofpacket
	wire   [90:0] cmd_xbar_demux_002_src1_data;                                                                                                     // cmd_xbar_demux_002:src1_data -> width_adapter_005:in_data
	wire   [18:0] cmd_xbar_demux_002_src1_channel;                                                                                                  // cmd_xbar_demux_002:src1_channel -> width_adapter_005:in_channel
	wire          cmd_xbar_demux_002_src1_ready;                                                                                                    // width_adapter_005:in_ready -> cmd_xbar_demux_002:src1_ready
	wire          width_adapter_005_src_endofpacket;                                                                                                // width_adapter_005:out_endofpacket -> cmd_xbar_mux_018:sink1_endofpacket
	wire          width_adapter_005_src_valid;                                                                                                      // width_adapter_005:out_valid -> cmd_xbar_mux_018:sink1_valid
	wire          width_adapter_005_src_startofpacket;                                                                                              // width_adapter_005:out_startofpacket -> cmd_xbar_mux_018:sink1_startofpacket
	wire  [108:0] width_adapter_005_src_data;                                                                                                       // width_adapter_005:out_data -> cmd_xbar_mux_018:sink1_data
	wire          width_adapter_005_src_ready;                                                                                                      // cmd_xbar_mux_018:sink1_ready -> width_adapter_005:out_ready
	wire   [18:0] width_adapter_005_src_channel;                                                                                                    // width_adapter_005:out_channel -> cmd_xbar_mux_018:sink1_channel
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                                              // rsp_xbar_demux_002:src0_endofpacket -> width_adapter_006:in_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                                                    // rsp_xbar_demux_002:src0_valid -> width_adapter_006:in_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                                                            // rsp_xbar_demux_002:src0_startofpacket -> width_adapter_006:in_startofpacket
	wire   [90:0] rsp_xbar_demux_002_src0_data;                                                                                                     // rsp_xbar_demux_002:src0_data -> width_adapter_006:in_data
	wire   [18:0] rsp_xbar_demux_002_src0_channel;                                                                                                  // rsp_xbar_demux_002:src0_channel -> width_adapter_006:in_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                                                    // width_adapter_006:in_ready -> rsp_xbar_demux_002:src0_ready
	wire          width_adapter_006_src_endofpacket;                                                                                                // width_adapter_006:out_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          width_adapter_006_src_valid;                                                                                                      // width_adapter_006:out_valid -> rsp_xbar_mux:sink2_valid
	wire          width_adapter_006_src_startofpacket;                                                                                              // width_adapter_006:out_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [108:0] width_adapter_006_src_data;                                                                                                       // width_adapter_006:out_data -> rsp_xbar_mux:sink2_data
	wire          width_adapter_006_src_ready;                                                                                                      // rsp_xbar_mux:sink2_ready -> width_adapter_006:out_ready
	wire   [18:0] width_adapter_006_src_channel;                                                                                                    // width_adapter_006:out_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src1_endofpacket;                                                                                              // rsp_xbar_demux_002:src1_endofpacket -> width_adapter_007:in_endofpacket
	wire          rsp_xbar_demux_002_src1_valid;                                                                                                    // rsp_xbar_demux_002:src1_valid -> width_adapter_007:in_valid
	wire          rsp_xbar_demux_002_src1_startofpacket;                                                                                            // rsp_xbar_demux_002:src1_startofpacket -> width_adapter_007:in_startofpacket
	wire   [90:0] rsp_xbar_demux_002_src1_data;                                                                                                     // rsp_xbar_demux_002:src1_data -> width_adapter_007:in_data
	wire   [18:0] rsp_xbar_demux_002_src1_channel;                                                                                                  // rsp_xbar_demux_002:src1_channel -> width_adapter_007:in_channel
	wire          rsp_xbar_demux_002_src1_ready;                                                                                                    // width_adapter_007:in_ready -> rsp_xbar_demux_002:src1_ready
	wire          width_adapter_007_src_endofpacket;                                                                                                // width_adapter_007:out_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          width_adapter_007_src_valid;                                                                                                      // width_adapter_007:out_valid -> rsp_xbar_mux_001:sink2_valid
	wire          width_adapter_007_src_startofpacket;                                                                                              // width_adapter_007:out_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [108:0] width_adapter_007_src_data;                                                                                                       // width_adapter_007:out_data -> rsp_xbar_mux_001:sink2_data
	wire          width_adapter_007_src_ready;                                                                                                      // rsp_xbar_mux_001:sink2_ready -> width_adapter_007:out_ready
	wire   [18:0] width_adapter_007_src_channel;                                                                                                    // width_adapter_007:out_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                                                              // rsp_xbar_demux_011:src0_endofpacket -> width_adapter_008:in_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                                                    // rsp_xbar_demux_011:src0_valid -> width_adapter_008:in_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                                                            // rsp_xbar_demux_011:src0_startofpacket -> width_adapter_008:in_startofpacket
	wire   [81:0] rsp_xbar_demux_011_src0_data;                                                                                                     // rsp_xbar_demux_011:src0_data -> width_adapter_008:in_data
	wire   [18:0] rsp_xbar_demux_011_src0_channel;                                                                                                  // rsp_xbar_demux_011:src0_channel -> width_adapter_008:in_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                                                    // width_adapter_008:in_ready -> rsp_xbar_demux_011:src0_ready
	wire          width_adapter_008_src_endofpacket;                                                                                                // width_adapter_008:out_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire          width_adapter_008_src_valid;                                                                                                      // width_adapter_008:out_valid -> rsp_xbar_mux_001:sink11_valid
	wire          width_adapter_008_src_startofpacket;                                                                                              // width_adapter_008:out_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [108:0] width_adapter_008_src_data;                                                                                                       // width_adapter_008:out_data -> rsp_xbar_mux_001:sink11_data
	wire          width_adapter_008_src_ready;                                                                                                      // rsp_xbar_mux_001:sink11_ready -> width_adapter_008:out_ready
	wire   [18:0] width_adapter_008_src_channel;                                                                                                    // width_adapter_008:out_channel -> rsp_xbar_mux_001:sink11_channel
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                                                              // rsp_xbar_demux_015:src0_endofpacket -> width_adapter_009:in_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                                                    // rsp_xbar_demux_015:src0_valid -> width_adapter_009:in_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                                                            // rsp_xbar_demux_015:src0_startofpacket -> width_adapter_009:in_startofpacket
	wire   [81:0] rsp_xbar_demux_015_src0_data;                                                                                                     // rsp_xbar_demux_015:src0_data -> width_adapter_009:in_data
	wire   [18:0] rsp_xbar_demux_015_src0_channel;                                                                                                  // rsp_xbar_demux_015:src0_channel -> width_adapter_009:in_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                                                    // width_adapter_009:in_ready -> rsp_xbar_demux_015:src0_ready
	wire          width_adapter_009_src_endofpacket;                                                                                                // width_adapter_009:out_endofpacket -> rsp_xbar_mux_001:sink15_endofpacket
	wire          width_adapter_009_src_valid;                                                                                                      // width_adapter_009:out_valid -> rsp_xbar_mux_001:sink15_valid
	wire          width_adapter_009_src_startofpacket;                                                                                              // width_adapter_009:out_startofpacket -> rsp_xbar_mux_001:sink15_startofpacket
	wire  [108:0] width_adapter_009_src_data;                                                                                                       // width_adapter_009:out_data -> rsp_xbar_mux_001:sink15_data
	wire          width_adapter_009_src_ready;                                                                                                      // rsp_xbar_mux_001:sink15_ready -> width_adapter_009:out_ready
	wire   [18:0] width_adapter_009_src_channel;                                                                                                    // width_adapter_009:out_channel -> rsp_xbar_mux_001:sink15_channel
	wire          rsp_xbar_demux_016_src0_endofpacket;                                                                                              // rsp_xbar_demux_016:src0_endofpacket -> width_adapter_010:in_endofpacket
	wire          rsp_xbar_demux_016_src0_valid;                                                                                                    // rsp_xbar_demux_016:src0_valid -> width_adapter_010:in_valid
	wire          rsp_xbar_demux_016_src0_startofpacket;                                                                                            // rsp_xbar_demux_016:src0_startofpacket -> width_adapter_010:in_startofpacket
	wire   [90:0] rsp_xbar_demux_016_src0_data;                                                                                                     // rsp_xbar_demux_016:src0_data -> width_adapter_010:in_data
	wire   [18:0] rsp_xbar_demux_016_src0_channel;                                                                                                  // rsp_xbar_demux_016:src0_channel -> width_adapter_010:in_channel
	wire          rsp_xbar_demux_016_src0_ready;                                                                                                    // width_adapter_010:in_ready -> rsp_xbar_demux_016:src0_ready
	wire          width_adapter_010_src_endofpacket;                                                                                                // width_adapter_010:out_endofpacket -> rsp_xbar_mux_001:sink16_endofpacket
	wire          width_adapter_010_src_valid;                                                                                                      // width_adapter_010:out_valid -> rsp_xbar_mux_001:sink16_valid
	wire          width_adapter_010_src_startofpacket;                                                                                              // width_adapter_010:out_startofpacket -> rsp_xbar_mux_001:sink16_startofpacket
	wire  [108:0] width_adapter_010_src_data;                                                                                                       // width_adapter_010:out_data -> rsp_xbar_mux_001:sink16_data
	wire          width_adapter_010_src_ready;                                                                                                      // rsp_xbar_mux_001:sink16_ready -> width_adapter_010:out_ready
	wire   [18:0] width_adapter_010_src_channel;                                                                                                    // width_adapter_010:out_channel -> rsp_xbar_mux_001:sink16_channel
	wire          rsp_xbar_demux_018_src1_endofpacket;                                                                                              // rsp_xbar_demux_018:src1_endofpacket -> width_adapter_011:in_endofpacket
	wire          rsp_xbar_demux_018_src1_valid;                                                                                                    // rsp_xbar_demux_018:src1_valid -> width_adapter_011:in_valid
	wire          rsp_xbar_demux_018_src1_startofpacket;                                                                                            // rsp_xbar_demux_018:src1_startofpacket -> width_adapter_011:in_startofpacket
	wire  [108:0] rsp_xbar_demux_018_src1_data;                                                                                                     // rsp_xbar_demux_018:src1_data -> width_adapter_011:in_data
	wire   [18:0] rsp_xbar_demux_018_src1_channel;                                                                                                  // rsp_xbar_demux_018:src1_channel -> width_adapter_011:in_channel
	wire          rsp_xbar_demux_018_src1_ready;                                                                                                    // width_adapter_011:in_ready -> rsp_xbar_demux_018:src1_ready
	wire          width_adapter_011_src_endofpacket;                                                                                                // width_adapter_011:out_endofpacket -> rsp_xbar_mux_002:sink1_endofpacket
	wire          width_adapter_011_src_valid;                                                                                                      // width_adapter_011:out_valid -> rsp_xbar_mux_002:sink1_valid
	wire          width_adapter_011_src_startofpacket;                                                                                              // width_adapter_011:out_startofpacket -> rsp_xbar_mux_002:sink1_startofpacket
	wire   [90:0] width_adapter_011_src_data;                                                                                                       // width_adapter_011:out_data -> rsp_xbar_mux_002:sink1_data
	wire          width_adapter_011_src_ready;                                                                                                      // rsp_xbar_mux_002:sink1_ready -> width_adapter_011:out_ready
	wire   [18:0] width_adapter_011_src_channel;                                                                                                    // width_adapter_011:out_channel -> rsp_xbar_mux_002:sink1_channel
	wire   [18:0] limiter_cmd_valid_data;                                                                                                           // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire   [18:0] limiter_001_cmd_valid_data;                                                                                                       // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	wire   [18:0] limiter_002_cmd_valid_data;                                                                                                       // limiter_002:cmd_src_valid -> cmd_xbar_demux_002:sink_valid
	wire          irq_mapper_receiver0_irq;                                                                                                         // JTAG:av_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                                                                         // sdcard_timer:irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                                                                                         // ps2_0:irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                                                                                         // audio_0:irq -> irq_mapper:receiver3_irq
	wire          irq_mapper_receiver4_irq;                                                                                                         // usb_0:irq -> irq_mapper:receiver4_irq
	wire   [31:0] nios2_system_d_irq_irq;                                                                                                           // irq_mapper:sender_irq -> nios2_system:d_irq

	nios2_system_nios2_system nios2_system (
		.clk                                   (clocks_sys_clk_clk),                                                        //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                           //                   reset_n.reset_n
		.d_address                             (nios2_system_data_master_address),                                          //               data_master.address
		.d_byteenable                          (nios2_system_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (nios2_system_data_master_read),                                             //                          .read
		.d_readdata                            (nios2_system_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (nios2_system_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (nios2_system_data_master_write),                                            //                          .write
		.d_writedata                           (nios2_system_data_master_writedata),                                        //                          .writedata
		.d_readdatavalid                       (nios2_system_data_master_readdatavalid),                                    //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_system_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (nios2_system_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (nios2_system_instruction_master_read),                                      //                          .read
		.i_readdata                            (nios2_system_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (nios2_system_instruction_master_waitrequest),                               //                          .waitrequest
		.i_readdatavalid                       (nios2_system_instruction_master_readdatavalid),                             //                          .readdatavalid
		.d_irq                                 (nios2_system_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_system_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_system_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (nios2_system_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_system_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (nios2_system_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (nios2_system_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (nios2_system_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (nios2_system_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (nios2_system_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                           // custom_instruction_master.readra
	);

	nios2_system_clocks clocks (
		.CLOCK_50    (clk_clk),                            //       clk_in_primary.clk
		.reset       (rst_controller_001_reset_out_reset), // clk_in_primary_reset.reset
		.sys_clk     (clocks_sys_clk_clk),                 //              sys_clk.clk
		.sys_reset_n (),                                   //        sys_clk_reset.reset_n
		.SDRAM_CLK   (sdram_clk_clk),                      //            sdram_clk.clk
		.VGA_CLK     (clocks_vga_clk_clk),                 //              vga_clk.clk
		.CLOCK_27    (audio_secondary_clk),                //     clk_in_secondary.clk
		.AUD_CLK     (audio_clk_clk)                       //            audio_clk.clk
	);

	nios2_system_onchip onchip (
		.clk        (clocks_sys_clk_clk),                                  //   clk1.clk
		.address    (onchip_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (onchip_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (onchip_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (onchip_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (onchip_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (onchip_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                   //       .reset_req
	);

	nios2_system_sdram sdram (
		.clk            (clocks_sys_clk_clk),                                    //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                       // reset.reset_n
		.az_addr        (sdram_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                                       //  wire.export
		.zs_ba          (sdram_wire_ba),                                         //      .export
		.zs_cas_n       (sdram_wire_cas_n),                                      //      .export
		.zs_cke         (sdram_wire_cke),                                        //      .export
		.zs_cs_n        (sdram_wire_cs_n),                                       //      .export
		.zs_dq          (sdram_wire_dq),                                         //      .export
		.zs_dqm         (sdram_wire_dqm),                                        //      .export
		.zs_ras_n       (sdram_wire_ras_n),                                      //      .export
		.zs_we_n        (sdram_wire_we_n)                                        //      .export
	);

	nios2_system_LEDG ledg (
		.clk        (clocks_sys_clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (ledg_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ledg_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ledg_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ledg_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ledg_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ledg_export)                                        // external_connection.export
	);

	nios2_system_LEDR ledr (
		.clk        (clocks_sys_clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (ledr_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ledr_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ledr_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ledr_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ledr_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ledr_export)                                        // external_connection.export
	);

	nios2_system_switches switches (
		.clk      (clocks_sys_clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address  (switches_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (switches_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (switches_export)                                      // external_connection.export
	);

	nios2_system_key key (
		.clk      (clocks_sys_clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (key_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (key_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (keys_export)                                     // external_connection.export
	);

	nios2_system_character_lcd_0 character_lcd_0 (
		.clk         (clocks_sys_clk_clk),                                                          //        clock_reset.clk
		.reset       (rst_controller_reset_out_reset),                                              //  clock_reset_reset.reset
		.address     (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_address),     //   avalon_lcd_slave.address
		.chipselect  (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_chipselect),  //                   .chipselect
		.read        (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_read),        //                   .read
		.write       (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_write),       //                   .write
		.writedata   (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_writedata),   //                   .writedata
		.readdata    (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_readdata),    //                   .readdata
		.waitrequest (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_waitrequest), //                   .waitrequest
		.LCD_DATA    (lcd_data_DATA),                                                               // external_interface.export
		.LCD_ON      (lcd_data_ON),                                                                 //                   .export
		.LCD_BLON    (lcd_data_BLON),                                                               //                   .export
		.LCD_EN      (lcd_data_EN),                                                                 //                   .export
		.LCD_RS      (lcd_data_RS),                                                                 //                   .export
		.LCD_RW      (lcd_data_RW)                                                                  //                   .export
	);

	nios2_system_JTAG jtag (
		.clk            (clocks_sys_clk_clk),                                                //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                   //             reset.reset_n
		.av_chipselect  (jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                           //               irq.irq
	);

	nios2_system_video_pixel_buffer_dma video_pixel_buffer_dma (
		.clk                  (clocks_sys_clk_clk),                                                                    //             clock_reset.clk
		.reset                (rst_controller_reset_out_reset),                                                        //       clock_reset_reset.reset
		.master_readdatavalid (video_pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid),                          // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (video_pixel_buffer_dma_avalon_pixel_dma_master_waitrequest),                            //                        .waitrequest
		.master_address       (video_pixel_buffer_dma_avalon_pixel_dma_master_address),                                //                        .address
		.master_arbiterlock   (video_pixel_buffer_dma_avalon_pixel_dma_master_lock),                                   //                        .lock
		.master_read          (video_pixel_buffer_dma_avalon_pixel_dma_master_read),                                   //                        .read
		.master_readdata      (video_pixel_buffer_dma_avalon_pixel_dma_master_readdata),                               //                        .readdata
		.slave_address        (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_address),    //    avalon_control_slave.address
		.slave_byteenable     (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_byteenable), //                        .byteenable
		.slave_read           (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_read),       //                        .read
		.slave_write          (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_write),      //                        .write
		.slave_writedata      (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_writedata),  //                        .writedata
		.slave_readdata       (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_readdata),   //                        .readdata
		.stream_ready         (video_pixel_buffer_dma_avalon_pixel_source_ready),                                      //     avalon_pixel_source.ready
		.stream_startofpacket (video_pixel_buffer_dma_avalon_pixel_source_startofpacket),                              //                        .startofpacket
		.stream_endofpacket   (video_pixel_buffer_dma_avalon_pixel_source_endofpacket),                                //                        .endofpacket
		.stream_valid         (video_pixel_buffer_dma_avalon_pixel_source_valid),                                      //                        .valid
		.stream_data          (video_pixel_buffer_dma_avalon_pixel_source_data)                                        //                        .data
	);

	nios2_system_video_rgb_resampler_0 video_rgb_resampler_0 (
		.clk                      (clocks_sys_clk_clk),                                       //       clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                           // clock_reset_reset.reset
		.stream_in_startofpacket  (video_pixel_buffer_dma_avalon_pixel_source_startofpacket), //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (video_pixel_buffer_dma_avalon_pixel_source_endofpacket),   //                  .endofpacket
		.stream_in_valid          (video_pixel_buffer_dma_avalon_pixel_source_valid),         //                  .valid
		.stream_in_ready          (video_pixel_buffer_dma_avalon_pixel_source_ready),         //                  .ready
		.stream_in_data           (video_pixel_buffer_dma_avalon_pixel_source_data),          //                  .data
		.stream_out_ready         (video_rgb_resampler_0_avalon_rgb_source_ready),            // avalon_rgb_source.ready
		.stream_out_startofpacket (video_rgb_resampler_0_avalon_rgb_source_startofpacket),    //                  .startofpacket
		.stream_out_endofpacket   (video_rgb_resampler_0_avalon_rgb_source_endofpacket),      //                  .endofpacket
		.stream_out_valid         (video_rgb_resampler_0_avalon_rgb_source_valid),            //                  .valid
		.stream_out_data          (video_rgb_resampler_0_avalon_rgb_source_data)              //                  .data
	);

	nios2_system_video_scaler_0 video_scaler_0 (
		.clk                      (clocks_sys_clk_clk),                                    //          clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                        //    clock_reset_reset.reset
		.stream_in_startofpacket  (video_rgb_resampler_0_avalon_rgb_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (video_rgb_resampler_0_avalon_rgb_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (video_rgb_resampler_0_avalon_rgb_source_valid),         //                     .valid
		.stream_in_ready          (video_rgb_resampler_0_avalon_rgb_source_ready),         //                     .ready
		.stream_in_data           (video_rgb_resampler_0_avalon_rgb_source_data),          //                     .data
		.stream_out_ready         (video_scaler_0_avalon_scaler_source_ready),             // avalon_scaler_source.ready
		.stream_out_startofpacket (video_scaler_0_avalon_scaler_source_startofpacket),     //                     .startofpacket
		.stream_out_endofpacket   (video_scaler_0_avalon_scaler_source_endofpacket),       //                     .endofpacket
		.stream_out_valid         (video_scaler_0_avalon_scaler_source_valid),             //                     .valid
		.stream_out_data          (video_scaler_0_avalon_scaler_source_data)               //                     .data
	);

	nios2_system_video_dual_clock_buffer_0 video_dual_clock_buffer_0 (
		.clk_stream_in            (clocks_sys_clk_clk),                                              //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_reset_out_reset),                                  //   clock_stream_in_reset.reset
		.clk_stream_out           (clocks_vga_clk_clk),                                              //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_002_reset_out_reset),                              //  clock_stream_out_reset.reset
		.stream_in_ready          (video_alpha_blender_0_avalon_blended_source_ready),               //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (video_alpha_blender_0_avalon_blended_source_startofpacket),       //                        .startofpacket
		.stream_in_endofpacket    (video_alpha_blender_0_avalon_blended_source_endofpacket),         //                        .endofpacket
		.stream_in_valid          (video_alpha_blender_0_avalon_blended_source_valid),               //                        .valid
		.stream_in_data           (video_alpha_blender_0_avalon_blended_source_data),                //                        .data
		.stream_out_ready         (video_dual_clock_buffer_0_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (video_dual_clock_buffer_0_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (video_dual_clock_buffer_0_avalon_dc_buffer_source_data)           //                        .data
	);

	nios2_system_video_vga_controller_0 video_vga_controller_0 (
		.clk           (clocks_vga_clk_clk),                                              //        clock_reset.clk
		.reset         (rst_controller_002_reset_out_reset),                              //  clock_reset_reset.reset
		.data          (video_dual_clock_buffer_0_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (video_dual_clock_buffer_0_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (video_dual_clock_buffer_0_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (video_vga_controller_0_external_interface_CLK),                   // external_interface.export
		.VGA_HS        (video_vga_controller_0_external_interface_HS),                    //                   .export
		.VGA_VS        (video_vga_controller_0_external_interface_VS),                    //                   .export
		.VGA_BLANK     (video_vga_controller_0_external_interface_BLANK),                 //                   .export
		.VGA_SYNC      (video_vga_controller_0_external_interface_SYNC),                  //                   .export
		.VGA_R         (video_vga_controller_0_external_interface_R),                     //                   .export
		.VGA_G         (video_vga_controller_0_external_interface_G),                     //                   .export
		.VGA_B         (video_vga_controller_0_external_interface_B)                      //                   .export
	);

	nios2_system_video_character_buffer_with_dma_0 video_character_buffer_with_dma_0 (
		.clk                  (clocks_sys_clk_clk),                                                                                    //               clock_reset.clk
		.reset                (rst_controller_reset_out_reset),                                                                        //         clock_reset_reset.reset
		.ctrl_address         (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_anti_slave_0_address),    // avalon_char_control_slave.address
		.ctrl_byteenable      (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_anti_slave_0_byteenable), //                          .byteenable
		.ctrl_chipselect      (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_anti_slave_0_chipselect), //                          .chipselect
		.ctrl_read            (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_anti_slave_0_read),       //                          .read
		.ctrl_write           (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_anti_slave_0_write),      //                          .write
		.ctrl_writedata       (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_anti_slave_0_writedata),  //                          .writedata
		.ctrl_readdata        (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_anti_slave_0_readdata),   //                          .readdata
		.buf_byteenable       (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_anti_slave_0_byteenable),  //  avalon_char_buffer_slave.byteenable
		.buf_chipselect       (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_anti_slave_0_chipselect),  //                          .chipselect
		.buf_read             (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_anti_slave_0_read),        //                          .read
		.buf_write            (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_anti_slave_0_write),       //                          .write
		.buf_writedata        (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.buf_readdata         (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.buf_waitrequest      (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.buf_address          (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_anti_slave_0_address),     //                          .address
		.stream_ready         (video_character_buffer_with_dma_0_avalon_char_source_ready),                                            //        avalon_char_source.ready
		.stream_startofpacket (video_character_buffer_with_dma_0_avalon_char_source_startofpacket),                                    //                          .startofpacket
		.stream_endofpacket   (video_character_buffer_with_dma_0_avalon_char_source_endofpacket),                                      //                          .endofpacket
		.stream_valid         (video_character_buffer_with_dma_0_avalon_char_source_valid),                                            //                          .valid
		.stream_data          (video_character_buffer_with_dma_0_avalon_char_source_data)                                              //                          .data
	);

	nios2_system_video_alpha_blender_0 video_alpha_blender_0 (
		.clk                      (clocks_sys_clk_clk),                                                 //            clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                                     //      clock_reset_reset.reset
		.foreground_data          (video_character_buffer_with_dma_0_avalon_char_source_data),          // avalon_foreground_sink.data
		.foreground_startofpacket (video_character_buffer_with_dma_0_avalon_char_source_startofpacket), //                       .startofpacket
		.foreground_endofpacket   (video_character_buffer_with_dma_0_avalon_char_source_endofpacket),   //                       .endofpacket
		.foreground_valid         (video_character_buffer_with_dma_0_avalon_char_source_valid),         //                       .valid
		.foreground_ready         (video_character_buffer_with_dma_0_avalon_char_source_ready),         //                       .ready
		.background_data          (video_scaler_0_avalon_scaler_source_data),                           // avalon_background_sink.data
		.background_startofpacket (video_scaler_0_avalon_scaler_source_startofpacket),                  //                       .startofpacket
		.background_endofpacket   (video_scaler_0_avalon_scaler_source_endofpacket),                    //                       .endofpacket
		.background_valid         (video_scaler_0_avalon_scaler_source_valid),                          //                       .valid
		.background_ready         (video_scaler_0_avalon_scaler_source_ready),                          //                       .ready
		.output_ready             (video_alpha_blender_0_avalon_blended_source_ready),                  //  avalon_blended_source.ready
		.output_data              (video_alpha_blender_0_avalon_blended_source_data),                   //                       .data
		.output_startofpacket     (video_alpha_blender_0_avalon_blended_source_startofpacket),          //                       .startofpacket
		.output_endofpacket       (video_alpha_blender_0_avalon_blended_source_endofpacket),            //                       .endofpacket
		.output_valid             (video_alpha_blender_0_avalon_blended_source_valid)                   //                       .valid
	);

	nios2_system_sdcard_timer sdcard_timer (
		.clk        (clocks_sys_clk_clk),                                        //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                           // reset.reset_n
		.address    (sdcard_timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (sdcard_timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (sdcard_timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (sdcard_timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~sdcard_timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                                   //   irq.irq
	);

	Altera_UP_SD_Card_Avalon_Interface altera_up_sd_card_avalon_interface_0 (
		.i_avalon_chip_select (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_sdcard_slave.chipselect
		.i_avalon_address     (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_address),     //                    .address
		.i_avalon_read        (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_read),        //                    .read
		.i_avalon_write       (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_write),       //                    .write
		.i_avalon_byteenable  (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_byteenable),  //                    .byteenable
		.i_avalon_writedata   (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_writedata),   //                    .writedata
		.o_avalon_readdata    (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_readdata),    //                    .readdata
		.o_avalon_waitrequest (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_waitrequest), //                    .waitrequest
		.i_clock              (clocks_sys_clk_clk),                                                                                  //          clock_sink.clk
		.i_reset_n            (~rst_controller_reset_out_reset),                                                                     //    clock_sink_reset.reset_n
		.b_SD_cmd             (sdcard_b_SD_cmd),                                                                                     //         conduit_end.export
		.b_SD_dat             (sdcard_b_SD_dat),                                                                                     //                    .export
		.b_SD_dat3            (sdcard_b_SD_dat3),                                                                                    //                    .export
		.o_SD_clock           (sdcard_o_SD_clock)                                                                                    //                    .export
	);

	nios2_system_ps2_0 ps2_0 (
		.clk         (clocks_sys_clk_clk),                                                //        clock_reset.clk
		.reset       (rst_controller_reset_out_reset),                                    //  clock_reset_reset.reset
		.address     (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_address),     //   avalon_ps2_slave.address
		.chipselect  (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_chipselect),  //                   .chipselect
		.byteenable  (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_byteenable),  //                   .byteenable
		.read        (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_read),        //                   .read
		.write       (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_write),       //                   .write
		.writedata   (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_writedata),   //                   .writedata
		.readdata    (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_readdata),    //                   .readdata
		.waitrequest (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_waitrequest), //                   .waitrequest
		.irq         (irq_mapper_receiver2_irq),                                          //          interrupt.irq
		.PS2_CLK     (ps2_peri_CLK),                                                      // external_interface.export
		.PS2_DAT     (ps2_peri_DAT)                                                       //                   .export
	);

	nios2_system_sram_0 sram_0 (
		.clk           (clocks_sys_clk_clk),                                                    //        clock_reset.clk
		.reset         (rst_controller_reset_out_reset),                                        //  clock_reset_reset.reset
		.SRAM_DQ       (sram_0_external_interface_DQ),                                          // external_interface.export
		.SRAM_ADDR     (sram_0_external_interface_ADDR),                                        //                   .export
		.SRAM_LB_N     (sram_0_external_interface_LB_N),                                        //                   .export
		.SRAM_UB_N     (sram_0_external_interface_UB_N),                                        //                   .export
		.SRAM_CE_N     (sram_0_external_interface_CE_N),                                        //                   .export
		.SRAM_OE_N     (sram_0_external_interface_OE_N),                                        //                   .export
		.SRAM_WE_N     (sram_0_external_interface_WE_N),                                        //                   .export
		.address       (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_address),       //  avalon_sram_slave.address
		.byteenable    (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),    //                   .byteenable
		.read          (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_read),          //                   .read
		.write         (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_write),         //                   .write
		.writedata     (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),     //                   .writedata
		.readdata      (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),      //                   .readdata
		.readdatavalid (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid)  //                   .readdatavalid
	);

	nios2_system_audio_0 audio_0 (
		.clk         (clocks_sys_clk_clk),                                                   //        clock_reset.clk
		.reset       (rst_controller_reset_out_reset),                                       //  clock_reset_reset.reset
		.address     (audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_address),    // avalon_audio_slave.address
		.chipselect  (audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_chipselect), //                   .chipselect
		.read        (audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_read),       //                   .read
		.write       (audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_write),      //                   .write
		.writedata   (audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_writedata),  //                   .writedata
		.readdata    (audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_readdata),   //                   .readdata
		.irq         (irq_mapper_receiver3_irq),                                             //          interrupt.irq
		.AUD_ADCDAT  (audio_ADCDAT),                                                         // external_interface.export
		.AUD_ADCLRCK (audio_ADCLRCK),                                                        //                   .export
		.AUD_BCLK    (audio_BCLK),                                                           //                   .export
		.AUD_DACDAT  (audio_DACDAT),                                                         //                   .export
		.AUD_DACLRCK (audio_DACLRCK)                                                         //                   .export
	);

	nios2_system_audio_and_video_config_0 audio_and_video_config_0 (
		.clk         (clocks_sys_clk_clk),                                                                         //            clock_reset.clk
		.reset       (rst_controller_reset_out_reset),                                                             //      clock_reset_reset.reset
		.address     (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_address),     // avalon_av_config_slave.address
		.byteenable  (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable),  //                       .byteenable
		.read        (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_read),        //                       .read
		.write       (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_write),       //                       .write
		.writedata   (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata),   //                       .writedata
		.readdata    (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata),    //                       .readdata
		.waitrequest (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest), //                       .waitrequest
		.I2C_SDAT    (av_config_SDAT),                                                                             //     external_interface.export
		.I2C_SCLK    (av_config_SCLK)                                                                              //                       .export
	);

	nios2_system_usb_0 usb_0 (
		.clk        (clocks_sys_clk_clk),                                               //        clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                                   //  clock_reset_reset.reset
		.address    (usb_0_avalon_usb_slave_translator_avalon_anti_slave_0_address),    //   avalon_usb_slave.address
		.chipselect (usb_0_avalon_usb_slave_translator_avalon_anti_slave_0_chipselect), //                   .chipselect
		.read       (usb_0_avalon_usb_slave_translator_avalon_anti_slave_0_read),       //                   .read
		.write      (usb_0_avalon_usb_slave_translator_avalon_anti_slave_0_write),      //                   .write
		.writedata  (usb_0_avalon_usb_slave_translator_avalon_anti_slave_0_writedata),  //                   .writedata
		.readdata   (usb_0_avalon_usb_slave_translator_avalon_anti_slave_0_readdata),   //                   .readdata
		.irq        (irq_mapper_receiver4_irq),                                         //          interrupt.irq
		.OTG_INT1   (usb_INT1),                                                         // external_interface.export
		.OTG_DATA   (usb_DATA),                                                         //                   .export
		.OTG_RST_N  (usb_RST_N),                                                        //                   .export
		.OTG_ADDR   (usb_ADDR),                                                         //                   .export
		.OTG_CS_N   (usb_CS_N),                                                         //                   .export
		.OTG_RD_N   (usb_RD_N),                                                         //                   .export
		.OTG_WR_N   (usb_WR_N),                                                         //                   .export
		.OTG_INT0   (usb_INT0)                                                          //                   .export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_system_instruction_master_translator (
		.clk                      (clocks_sys_clk_clk),                                                                 //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                     //                     reset.reset
		.uav_address              (nios2_system_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_system_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_system_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_system_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_system_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_system_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_system_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_system_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_system_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_system_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_system_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_system_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_system_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (nios2_system_instruction_master_read),                                               //                          .read
		.av_readdata              (nios2_system_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (nios2_system_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount            (1'b1),                                                                               //               (terminated)
		.av_byteenable            (4'b1111),                                                                            //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                               //               (terminated)
		.av_begintransfer         (1'b0),                                                                               //               (terminated)
		.av_chipselect            (1'b0),                                                                               //               (terminated)
		.av_write                 (1'b0),                                                                               //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                               //               (terminated)
		.av_lock                  (1'b0),                                                                               //               (terminated)
		.av_debugaccess           (1'b0),                                                                               //               (terminated)
		.uav_clken                (),                                                                                   //               (terminated)
		.av_clken                 (1'b1),                                                                               //               (terminated)
		.uav_response             (2'b00),                                                                              //               (terminated)
		.av_response              (),                                                                                   //               (terminated)
		.uav_writeresponserequest (),                                                                                   //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                               //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                               //               (terminated)
		.av_writeresponsevalid    ()                                                                                    //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_system_data_master_translator (
		.clk                      (clocks_sys_clk_clk),                                                          //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address              (nios2_system_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_system_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_system_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_system_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_system_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_system_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_system_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_system_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_system_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_system_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_system_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_system_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_system_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (nios2_system_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (nios2_system_data_master_read),                                               //                          .read
		.av_readdata              (nios2_system_data_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (nios2_system_data_master_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (nios2_system_data_master_write),                                              //                          .write
		.av_writedata             (nios2_system_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (nios2_system_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                                        //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                        //               (terminated)
		.av_begintransfer         (1'b0),                                                                        //               (terminated)
		.av_chipselect            (1'b0),                                                                        //               (terminated)
		.av_lock                  (1'b0),                                                                        //               (terminated)
		.uav_clken                (),                                                                            //               (terminated)
		.av_clken                 (1'b1),                                                                        //               (terminated)
		.uav_response             (2'b00),                                                                       //               (terminated)
		.av_response              (),                                                                            //               (terminated)
		.uav_writeresponserequest (),                                                                            //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                        //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                        //               (terminated)
		.av_writeresponsevalid    ()                                                                             //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) video_pixel_buffer_dma_avalon_pixel_dma_master_translator (
		.clk                      (clocks_sys_clk_clk),                                                                                //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                    //                     reset.reset
		.uav_address              (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (video_pixel_buffer_dma_avalon_pixel_dma_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (video_pixel_buffer_dma_avalon_pixel_dma_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (video_pixel_buffer_dma_avalon_pixel_dma_master_read),                                               //                          .read
		.av_readdata              (video_pixel_buffer_dma_avalon_pixel_dma_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (video_pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid),                                      //                          .readdatavalid
		.av_lock                  (video_pixel_buffer_dma_avalon_pixel_dma_master_lock),                                               //                          .lock
		.av_burstcount            (1'b1),                                                                                              //               (terminated)
		.av_byteenable            (2'b11),                                                                                             //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                                              //               (terminated)
		.av_begintransfer         (1'b0),                                                                                              //               (terminated)
		.av_chipselect            (1'b0),                                                                                              //               (terminated)
		.av_write                 (1'b0),                                                                                              //               (terminated)
		.av_writedata             (16'b0000000000000000),                                                                              //               (terminated)
		.av_debugaccess           (1'b0),                                                                                              //               (terminated)
		.uav_clken                (),                                                                                                  //               (terminated)
		.av_clken                 (1'b1),                                                                                              //               (terminated)
		.uav_response             (2'b00),                                                                                             //               (terminated)
		.av_response              (),                                                                                                  //               (terminated)
		.uav_writeresponserequest (),                                                                                                  //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                                              //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                                              //               (terminated)
		.av_writeresponsevalid    ()                                                                                                   //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_system_jtag_debug_module_translator (
		.clk                      (clocks_sys_clk_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                            //                    reset.reset
		.uav_address              (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (nios2_system_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (nios2_system_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (nios2_system_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (nios2_system_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (nios2_system_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (nios2_system_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (nios2_system_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (nios2_system_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                                          //              (terminated)
		.av_burstcount            (),                                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                                          //              (terminated)
		.av_lock                  (),                                                                                          //              (terminated)
		.av_chipselect            (),                                                                                          //              (terminated)
		.av_clken                 (),                                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                          //              (terminated)
		.uav_response             (),                                                                                          //              (terminated)
		.av_response              (2'b00),                                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_s1_translator (
		.clk                      (clocks_sys_clk_clk),                                                   //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address              (onchip_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (onchip_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (onchip_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (onchip_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (onchip_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (onchip_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (onchip_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (onchip_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (onchip_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (onchip_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (onchip_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (onchip_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (onchip_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (onchip_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (onchip_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (onchip_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (onchip_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (onchip_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                     //              (terminated)
		.av_begintransfer         (),                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                     //              (terminated)
		.av_burstcount            (),                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                     //              (terminated)
		.av_lock                  (),                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                 //              (terminated)
		.av_debugaccess           (),                                                                     //              (terminated)
		.av_outputenable          (),                                                                     //              (terminated)
		.uav_response             (),                                                                     //              (terminated)
		.av_response              (2'b00),                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_s1_translator (
		.clk                      (clocks_sys_clk_clk),                                                  //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sdram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sdram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sdram_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sdram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sdram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (sdram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (sdram_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (sdram_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (sdram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ledg_s1_translator (
		.clk                      (clocks_sys_clk_clk),                                                 //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (ledg_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ledg_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ledg_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ledg_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ledg_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ledg_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ledg_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ledg_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ledg_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ledg_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ledg_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ledg_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ledg_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ledg_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ledr_s1_translator (
		.clk                      (clocks_sys_clk_clk),                                                 //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (ledr_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ledr_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ledr_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ledr_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ledr_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ledr_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ledr_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ledr_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) switches_s1_translator (
		.clk                      (clocks_sys_clk_clk),                                                     //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                         //                    reset.reset
		.uav_address              (switches_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (switches_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (switches_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (switches_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (switches_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (switches_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (switches_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (switches_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (switches_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (switches_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (switches_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (switches_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (switches_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                       //              (terminated)
		.av_read                  (),                                                                       //              (terminated)
		.av_writedata             (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_chipselect            (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) key_s1_translator (
		.clk                      (clocks_sys_clk_clk),                                                //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                    //                    reset.reset
		.uav_address              (key_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (key_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (key_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (key_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (key_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (key_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (key_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (key_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (key_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (key_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (key_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (key_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (key_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                  //              (terminated)
		.av_read                  (),                                                                  //              (terminated)
		.av_writedata             (),                                                                  //              (terminated)
		.av_begintransfer         (),                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                  //              (terminated)
		.av_burstcount            (),                                                                  //              (terminated)
		.av_byteenable            (),                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                              //              (terminated)
		.av_writebyteenable       (),                                                                  //              (terminated)
		.av_lock                  (),                                                                  //              (terminated)
		.av_chipselect            (),                                                                  //              (terminated)
		.av_clken                 (),                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                              //              (terminated)
		.av_debugaccess           (),                                                                  //              (terminated)
		.av_outputenable          (),                                                                  //              (terminated)
		.uav_response             (),                                                                  //              (terminated)
		.av_response              (2'b00),                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdcard_timer_s1_translator (
		.clk                      (clocks_sys_clk_clk),                                                         //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                             //                    reset.reset
		.uav_address              (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sdcard_timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sdcard_timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (sdcard_timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sdcard_timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (sdcard_timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                           //              (terminated)
		.av_begintransfer         (),                                                                           //              (terminated)
		.av_beginbursttransfer    (),                                                                           //              (terminated)
		.av_burstcount            (),                                                                           //              (terminated)
		.av_byteenable            (),                                                                           //              (terminated)
		.av_readdatavalid         (1'b0),                                                                       //              (terminated)
		.av_waitrequest           (1'b0),                                                                       //              (terminated)
		.av_writebyteenable       (),                                                                           //              (terminated)
		.av_lock                  (),                                                                           //              (terminated)
		.av_clken                 (),                                                                           //              (terminated)
		.uav_clken                (1'b0),                                                                       //              (terminated)
		.av_debugaccess           (),                                                                           //              (terminated)
		.av_outputenable          (),                                                                           //              (terminated)
		.uav_response             (),                                                                           //              (terminated)
		.av_response              (2'b00),                                                                      //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                       //              (terminated)
		.uav_writeresponsevalid   (),                                                                           //              (terminated)
		.av_writeresponserequest  (),                                                                           //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (8),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator (
		.clk                      (clocks_sys_clk_clk),                                                                                                  //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                                      //                    reset.reset
		.uav_address              (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                                                                    //              (terminated)
		.av_burstcount            (),                                                                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                                                //              (terminated)
		.av_writebyteenable       (),                                                                                                                    //              (terminated)
		.av_lock                  (),                                                                                                                    //              (terminated)
		.av_clken                 (),                                                                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                                                                //              (terminated)
		.av_debugaccess           (),                                                                                                                    //              (terminated)
		.av_outputenable          (),                                                                                                                    //              (terminated)
		.uav_response             (),                                                                                                                    //              (terminated)
		.av_response              (2'b00),                                                                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ps2_0_avalon_ps2_slave_translator (
		.clk                      (clocks_sys_clk_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                    //                    reset.reset
		.uav_address              (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (ps2_0_avalon_ps2_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                                  //              (terminated)
		.av_burstcount            (),                                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                                              //              (terminated)
		.av_writebyteenable       (),                                                                                  //              (terminated)
		.av_lock                  (),                                                                                  //              (terminated)
		.av_clken                 (),                                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                                              //              (terminated)
		.av_debugaccess           (),                                                                                  //              (terminated)
		.av_outputenable          (),                                                                                  //              (terminated)
		.uav_response             (),                                                                                  //              (terminated)
		.av_response              (2'b00),                                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) audio_0_avalon_audio_slave_translator (
		.clk                      (clocks_sys_clk_clk),                                                                    //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                        //                    reset.reset
		.uav_address              (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (audio_0_avalon_audio_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                                      //              (terminated)
		.av_burstcount            (),                                                                                      //              (terminated)
		.av_byteenable            (),                                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                                      //              (terminated)
		.av_lock                  (),                                                                                      //              (terminated)
		.av_clken                 (),                                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                                  //              (terminated)
		.av_debugaccess           (),                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                      //              (terminated)
		.uav_response             (),                                                                                      //              (terminated)
		.av_response              (2'b00),                                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) character_lcd_0_avalon_lcd_slave_translator (
		.clk                      (clocks_sys_clk_clk),                                                                          //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                              //                    reset.reset
		.uav_address              (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                                            //              (terminated)
		.av_burstcount            (),                                                                                            //              (terminated)
		.av_byteenable            (),                                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                                            //              (terminated)
		.av_lock                  (),                                                                                            //              (terminated)
		.av_clken                 (),                                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                                        //              (terminated)
		.av_debugaccess           (),                                                                                            //              (terminated)
		.av_outputenable          (),                                                                                            //              (terminated)
		.uav_response             (),                                                                                            //              (terminated)
		.av_response              (2'b00),                                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_avalon_jtag_slave_translator (
		.clk                      (clocks_sys_clk_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                    //                    reset.reset
		.uav_address              (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                                  //              (terminated)
		.av_burstcount            (),                                                                                  //              (terminated)
		.av_byteenable            (),                                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                                              //              (terminated)
		.av_writebyteenable       (),                                                                                  //              (terminated)
		.av_lock                  (),                                                                                  //              (terminated)
		.av_clken                 (),                                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                                              //              (terminated)
		.av_debugaccess           (),                                                                                  //              (terminated)
		.av_outputenable          (),                                                                                  //              (terminated)
		.uav_response             (),                                                                                  //              (terminated)
		.av_response              (2'b00),                                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) video_pixel_buffer_dma_avalon_control_slave_translator (
		.clk                      (clocks_sys_clk_clk),                                                                                     //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                         //                    reset.reset
		.uav_address              (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_begintransfer         (),                                                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                                                       //              (terminated)
		.av_burstcount            (),                                                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                                                       //              (terminated)
		.av_lock                  (),                                                                                                       //              (terminated)
		.av_chipselect            (),                                                                                                       //              (terminated)
		.av_clken                 (),                                                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                                                   //              (terminated)
		.av_debugaccess           (),                                                                                                       //              (terminated)
		.av_outputenable          (),                                                                                                       //              (terminated)
		.uav_response             (),                                                                                                       //              (terminated)
		.av_response              (2'b00),                                                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) video_character_buffer_with_dma_0_avalon_char_control_slave_translator (
		.clk                      (clocks_sys_clk_clk),                                                                                                     //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                                         //                    reset.reset
		.uav_address              (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                                                                       //              (terminated)
		.av_burstcount            (),                                                                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                                                                       //              (terminated)
		.av_lock                  (),                                                                                                                       //              (terminated)
		.av_clken                 (),                                                                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                                                                   //              (terminated)
		.av_debugaccess           (),                                                                                                                       //              (terminated)
		.av_outputenable          (),                                                                                                                       //              (terminated)
		.uav_response             (),                                                                                                                       //              (terminated)
		.av_response              (2'b00),                                                                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (13),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator (
		.clk                      (clocks_sys_clk_clk),                                                                                                    //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                                        //                    reset.reset
		.uav_address              (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                                                                      //              (terminated)
		.av_burstcount            (),                                                                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                                                                      //              (terminated)
		.av_lock                  (),                                                                                                                      //              (terminated)
		.av_clken                 (),                                                                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                                                                  //              (terminated)
		.av_debugaccess           (),                                                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                                                      //              (terminated)
		.uav_response             (),                                                                                                                      //              (terminated)
		.av_response              (2'b00),                                                                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (18),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sram_0_avalon_sram_slave_translator (
		.clk                      (clocks_sys_clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                      //                    reset.reset
		.uav_address              (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_begintransfer         (),                                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                                    //              (terminated)
		.av_burstcount            (),                                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                                //              (terminated)
		.av_writebyteenable       (),                                                                                    //              (terminated)
		.av_lock                  (),                                                                                    //              (terminated)
		.av_chipselect            (),                                                                                    //              (terminated)
		.av_clken                 (),                                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                                //              (terminated)
		.av_debugaccess           (),                                                                                    //              (terminated)
		.av_outputenable          (),                                                                                    //              (terminated)
		.uav_response             (),                                                                                    //              (terminated)
		.av_response              (2'b00),                                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) audio_and_video_config_0_avalon_av_config_slave_translator (
		.clk                      (clocks_sys_clk_clk),                                                                                         //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                             //                    reset.reset
		.uav_address              (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer         (),                                                                                                           //              (terminated)
		.av_beginbursttransfer    (),                                                                                                           //              (terminated)
		.av_burstcount            (),                                                                                                           //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                                       //              (terminated)
		.av_writebyteenable       (),                                                                                                           //              (terminated)
		.av_lock                  (),                                                                                                           //              (terminated)
		.av_chipselect            (),                                                                                                           //              (terminated)
		.av_clken                 (),                                                                                                           //              (terminated)
		.uav_clken                (1'b0),                                                                                                       //              (terminated)
		.av_debugaccess           (),                                                                                                           //              (terminated)
		.av_outputenable          (),                                                                                                           //              (terminated)
		.uav_response             (),                                                                                                           //              (terminated)
		.av_response              (2'b00),                                                                                                      //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                                       //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                           //              (terminated)
		.av_writeresponserequest  (),                                                                                                           //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (5),
		.AV_WRITE_WAIT_CYCLES           (5),
		.AV_SETUP_WAIT_CYCLES           (5),
		.AV_DATA_HOLD_CYCLES            (5)
	) usb_0_avalon_usb_slave_translator (
		.clk                      (clocks_sys_clk_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                    //                    reset.reset
		.uav_address              (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (usb_0_avalon_usb_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (usb_0_avalon_usb_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (usb_0_avalon_usb_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (usb_0_avalon_usb_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (usb_0_avalon_usb_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (usb_0_avalon_usb_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                                  //              (terminated)
		.av_burstcount            (),                                                                                  //              (terminated)
		.av_byteenable            (),                                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                                              //              (terminated)
		.av_writebyteenable       (),                                                                                  //              (terminated)
		.av_lock                  (),                                                                                  //              (terminated)
		.av_clken                 (),                                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                                              //              (terminated)
		.av_debugaccess           (),                                                                                  //              (terminated)
		.av_outputenable          (),                                                                                  //              (terminated)
		.uav_response             (),                                                                                  //              (terminated)
		.av_response              (2'b00),                                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                               //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_THREAD_ID_H           (99),
		.PKT_THREAD_ID_L           (99),
		.PKT_CACHE_H               (106),
		.PKT_CACHE_L               (103),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.ST_DATA_W                 (109),
		.ST_CHANNEL_W              (19),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_system_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                          //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.av_address              (nios2_system_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_system_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_system_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_system_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_system_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_system_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_system_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_system_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_system_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_system_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_system_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_system_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_system_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_system_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_system_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_system_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_rsp_src_valid),                                                                       //        rp.valid
		.rp_data                 (limiter_rsp_src_data),                                                                        //          .data
		.rp_channel              (limiter_rsp_src_channel),                                                                     //          .channel
		.rp_startofpacket        (limiter_rsp_src_startofpacket),                                                               //          .startofpacket
		.rp_endofpacket          (limiter_rsp_src_endofpacket),                                                                 //          .endofpacket
		.rp_ready                (limiter_rsp_src_ready),                                                                       //          .ready
		.av_response             (),                                                                                            // (terminated)
		.av_writeresponserequest (1'b0),                                                                                        // (terminated)
		.av_writeresponsevalid   ()                                                                                             // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_THREAD_ID_H           (99),
		.PKT_THREAD_ID_L           (99),
		.PKT_CACHE_H               (106),
		.PKT_CACHE_L               (103),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.ST_DATA_W                 (109),
		.ST_CHANNEL_W              (19),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_system_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                   //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address              (nios2_system_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_system_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_system_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_system_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_system_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_system_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_system_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_system_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_system_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_system_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_system_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_system_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_system_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_system_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_system_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_system_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_001_rsp_src_valid),                                                            //        rp.valid
		.rp_data                 (limiter_001_rsp_src_data),                                                             //          .data
		.rp_channel              (limiter_001_rsp_src_channel),                                                          //          .channel
		.rp_startofpacket        (limiter_001_rsp_src_startofpacket),                                                    //          .startofpacket
		.rp_endofpacket          (limiter_001_rsp_src_endofpacket),                                                      //          .endofpacket
		.rp_ready                (limiter_001_rsp_src_ready),                                                            //          .ready
		.av_response             (),                                                                                     // (terminated)
		.av_writeresponserequest (1'b0),                                                                                 // (terminated)
		.av_writeresponsevalid   ()                                                                                      // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (76),
		.PKT_THREAD_ID_H           (81),
		.PKT_THREAD_ID_L           (81),
		.PKT_CACHE_H               (88),
		.PKT_CACHE_L               (85),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.ST_DATA_W                 (91),
		.ST_CHANNEL_W              (19),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (2),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                         //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                             // clk_reset.reset
		.av_address              (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_002_rsp_src_valid),                                                                                  //        rp.valid
		.rp_data                 (limiter_002_rsp_src_data),                                                                                   //          .data
		.rp_channel              (limiter_002_rsp_src_channel),                                                                                //          .channel
		.rp_startofpacket        (limiter_002_rsp_src_startofpacket),                                                                          //          .startofpacket
		.rp_endofpacket          (limiter_002_rsp_src_endofpacket),                                                                            //          .endofpacket
		.rp_ready                (limiter_002_rsp_src_ready),                                                                                  //          .ready
		.av_response             (),                                                                                                           // (terminated)
		.av_writeresponserequest (1'b0),                                                                                                       // (terminated)
		.av_writeresponsevalid   ()                                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                      //       clk_reset.reset
		.m0_address              (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                              //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                              //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                               //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                            //                .channel
		.rf_sink_ready           (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.in_data           (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) onchip_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (onchip_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                   //                .channel
		.rf_sink_ready           (onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (onchip_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (91),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                   //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                   //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                    //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                             //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                 //                .channel
		.rf_sink_ready           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (92),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (18),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clocks_sys_clk_clk),                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                   // (terminated)
		.csr_read          (1'b0),                                                                    // (terminated)
		.csr_write         (1'b0),                                                                    // (terminated)
		.csr_readdata      (),                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                    // (terminated)
		.almost_full_data  (),                                                                        // (terminated)
		.almost_empty_data (),                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                    // (terminated)
		.out_startofpacket (),                                                                        // (terminated)
		.out_endofpacket   (),                                                                        // (terminated)
		.in_empty          (1'b0),                                                                    // (terminated)
		.out_empty         (),                                                                        // (terminated)
		.in_error          (1'b0),                                                                    // (terminated)
		.out_error         (),                                                                        // (terminated)
		.in_channel        (1'b0),                                                                    // (terminated)
		.out_channel       ()                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ledg_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (ledg_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ledg_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ledg_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ledg_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ledg_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ledg_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ledg_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ledg_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ledg_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ledg_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ledg_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ledg_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ledg_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ledg_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_003_src_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_003_src_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_003_src_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_003_src_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_003_src_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_003_src_channel),                                                 //                .channel
		.rf_sink_ready           (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ledr_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (ledr_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ledr_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ledr_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ledr_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_004_src_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_004_src_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_004_src_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_004_src_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_004_src_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_004_src_channel),                                                 //                .channel
		.rf_sink_ready           (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) switches_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (switches_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (switches_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (switches_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (switches_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (switches_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (switches_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (switches_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (switches_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (switches_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (switches_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (switches_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (switches_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (switches_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (switches_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (switches_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (switches_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_005_src_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_mux_005_src_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_mux_005_src_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_mux_005_src_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_005_src_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_mux_005_src_channel),                                                     //                .channel
		.rf_sink_ready           (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) key_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (key_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (key_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (key_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (key_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (key_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (key_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (key_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (key_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (key_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (key_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (key_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (key_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (key_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (key_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (key_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (key_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_006_src_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_mux_006_src_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_mux_006_src_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_mux_006_src_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_006_src_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_mux_006_src_channel),                                                //                .channel
		.rf_sink_ready           (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (key_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (key_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (key_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (key_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (key_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.in_data           (key_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (key_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (key_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (key_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (key_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sdcard_timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_007_src_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_mux_007_src_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_mux_007_src_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_mux_007_src_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_007_src_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_mux_007_src_channel),                                                         //                .channel
		.rf_sink_ready           (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                //     (terminated)
		.m0_writeresponserequest (),                                                                                     //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                  //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                                //       clk_reset.reset
		.m0_address              (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_008_src_ready),                                                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_mux_008_src_valid),                                                                                                    //                .valid
		.cp_data                 (cmd_xbar_mux_008_src_data),                                                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_mux_008_src_startofpacket),                                                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_008_src_endofpacket),                                                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_mux_008_src_channel),                                                                                                  //                .channel
		.rf_sink_ready           (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                                                // clk_reset.reset
		.in_data           (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                                                          // (terminated)
		.csr_readdata      (),                                                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                                          // (terminated)
		.almost_full_data  (),                                                                                                                              // (terminated)
		.almost_empty_data (),                                                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                                                          // (terminated)
		.out_empty         (),                                                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                                                          // (terminated)
		.out_error         (),                                                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                                                          // (terminated)
		.out_channel       ()                                                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_009_src_ready),                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_mux_009_src_valid),                                                                  //                .valid
		.cp_data                 (cmd_xbar_mux_009_src_data),                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_mux_009_src_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_009_src_endofpacket),                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_mux_009_src_channel),                                                                //                .channel
		.rf_sink_ready           (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                  //       clk_reset.reset
		.m0_address              (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_010_src_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_010_src_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_010_src_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_010_src_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_010_src_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_010_src_channel),                                                                    //                .channel
		.rf_sink_ready           (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                  // clk_reset.reset
		.in_data           (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (60),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (66),
		.PKT_SRC_ID_L              (62),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (67),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (73),
		.PKT_RESPONSE_STATUS_H     (81),
		.PKT_RESPONSE_STATUS_L     (80),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                        //       clk_reset.reset
		.m0_address              (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                                       //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                                       //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                                        //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                                                     //                .channel
		.rf_sink_ready           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                        // clk_reset.reset
		.in_data           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                                  // (terminated)
		.csr_readdata      (),                                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                  // (terminated)
		.almost_full_data  (),                                                                                                      // (terminated)
		.almost_empty_data (),                                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                                  // (terminated)
		.out_empty         (),                                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                                  // (terminated)
		.out_error         (),                                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                                  // (terminated)
		.out_channel       ()                                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src12_ready),                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src12_valid),                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_001_src12_data),                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src12_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src12_endofpacket),                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src12_channel),                                                            //                .channel
		.rf_sink_ready           (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                   //       clk_reset.reset
		.m0_address              (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src13_ready),                                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src13_valid),                                                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src13_data),                                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src13_startofpacket),                                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src13_endofpacket),                                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src13_channel),                                                                                 //                .channel
		.rf_sink_ready           (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                                   // clk_reset.reset
		.in_data           (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                             // (terminated)
		.almost_full_data  (),                                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                                             // (terminated)
		.out_empty         (),                                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                                             // (terminated)
		.out_error         (),                                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                                             // (terminated)
		.out_channel       ()                                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                                   //       clk_reset.reset
		.m0_address              (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src14_ready),                                                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src14_valid),                                                                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src14_data),                                                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src14_startofpacket),                                                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src14_endofpacket),                                                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src14_channel),                                                                                                 //                .channel
		.rf_sink_ready           (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                                                   // clk_reset.reset
		.in_data           (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                                             // (terminated)
		.almost_full_data  (),                                                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                                                             // (terminated)
		.out_empty         (),                                                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                                                             // (terminated)
		.out_error         (),                                                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                                                             // (terminated)
		.out_channel       ()                                                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (60),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (66),
		.PKT_SRC_ID_L              (62),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (67),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (73),
		.PKT_RESPONSE_STATUS_H     (81),
		.PKT_RESPONSE_STATUS_L     (80),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                                  //       clk_reset.reset
		.m0_address              (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_002_source0_ready),                                                                                                 //              cp.ready
		.cp_valid                (burst_adapter_002_source0_valid),                                                                                                 //                .valid
		.cp_data                 (burst_adapter_002_source0_data),                                                                                                  //                .data
		.cp_startofpacket        (burst_adapter_002_source0_startofpacket),                                                                                         //                .startofpacket
		.cp_endofpacket          (burst_adapter_002_source0_endofpacket),                                                                                           //                .endofpacket
		.cp_channel              (burst_adapter_002_source0_channel),                                                                                               //                .channel
		.rf_sink_ready           (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                                                  // clk_reset.reset
		.in_data           (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                                            // (terminated)
		.almost_full_data  (),                                                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                                                            // (terminated)
		.out_empty         (),                                                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                                                            // (terminated)
		.out_error         (),                                                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                                                            // (terminated)
		.out_channel       ()                                                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (91),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                //       clk_reset.reset
		.m0_address              (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_003_source0_ready),                                                               //              cp.ready
		.cp_valid                (burst_adapter_003_source0_valid),                                                               //                .valid
		.cp_data                 (burst_adapter_003_source0_data),                                                                //                .data
		.cp_startofpacket        (burst_adapter_003_source0_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (burst_adapter_003_source0_endofpacket),                                                         //                .endofpacket
		.cp_channel              (burst_adapter_003_source0_channel),                                                             //                .channel
		.rf_sink_ready           (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (92),
		.FIFO_DEPTH          (3),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                // clk_reset.reset
		.in_data           (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (18),
		.FIFO_DEPTH          (3),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clocks_sys_clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                                    // (terminated)
		.out_startofpacket (),                                                                                        // (terminated)
		.out_endofpacket   (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                       //       clk_reset.reset
		.m0_address              (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src17_ready),                                                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src17_valid),                                                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_001_src17_data),                                                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src17_startofpacket),                                                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src17_endofpacket),                                                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src17_channel),                                                                                     //                .channel
		.rf_sink_ready           (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                                //     (terminated)
		.m0_writeresponserequest (),                                                                                                                     //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                                  //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                                       // clk_reset.reset
		.in_data           (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                                                 // (terminated)
		.csr_readdata      (),                                                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                                 // (terminated)
		.almost_full_data  (),                                                                                                                     // (terminated)
		.almost_empty_data (),                                                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                                                 // (terminated)
		.out_empty         (),                                                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                                                 // (terminated)
		.out_error         (),                                                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                                                 // (terminated)
		.out_channel       ()                                                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_018_src_ready),                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_mux_018_src_valid),                                                                  //                .valid
		.cp_data                 (cmd_xbar_mux_018_src_data),                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_mux_018_src_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_018_src_endofpacket),                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_mux_018_src_channel),                                                                //                .channel
		.rf_sink_ready           (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	nios2_system_addr_router addr_router (
		.sink_ready         (nios2_system_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_system_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_system_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_system_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_system_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                       //       src.ready
		.src_valid          (addr_router_src_valid),                                                                       //          .valid
		.src_data           (addr_router_src_data),                                                                        //          .data
		.src_channel        (addr_router_src_channel),                                                                     //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                               //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                                  //          .endofpacket
	);

	nios2_system_addr_router_001 addr_router_001 (
		.sink_ready         (nios2_system_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_system_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_system_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_system_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_system_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                            //          .valid
		.src_data           (addr_router_001_src_data),                                                             //          .data
		.src_channel        (addr_router_001_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                       //          .endofpacket
	);

	nios2_system_addr_router_002 addr_router_002 (
		.sink_ready         (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                             // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                                                  //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                                                  //          .valid
		.src_data           (addr_router_002_src_data),                                                                                   //          .data
		.src_channel        (addr_router_002_src_channel),                                                                                //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                                                          //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                                             //          .endofpacket
	);

	nios2_system_id_router id_router (
		.sink_ready         (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_system_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                       //       src.ready
		.src_valid          (id_router_src_valid),                                                                       //          .valid
		.src_data           (id_router_src_data),                                                                        //          .data
		.src_channel        (id_router_src_channel),                                                                     //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                               //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                                  //          .endofpacket
	);

	nios2_system_id_router id_router_001 (
		.sink_ready         (onchip_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                              //       src.ready
		.src_valid          (id_router_001_src_valid),                                              //          .valid
		.src_data           (id_router_001_src_data),                                               //          .data
		.src_channel        (id_router_001_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                         //          .endofpacket
	);

	nios2_system_id_router_002 id_router_002 (
		.sink_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                             //       src.ready
		.src_valid          (id_router_002_src_valid),                                             //          .valid
		.src_data           (id_router_002_src_data),                                              //          .data
		.src_channel        (id_router_002_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                        //          .endofpacket
	);

	nios2_system_id_router id_router_003 (
		.sink_ready         (ledg_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ledg_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ledg_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ledg_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ledg_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                            //       src.ready
		.src_valid          (id_router_003_src_valid),                                            //          .valid
		.src_data           (id_router_003_src_data),                                             //          .data
		.src_channel        (id_router_003_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                       //          .endofpacket
	);

	nios2_system_id_router id_router_004 (
		.sink_ready         (ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ledr_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                            //       src.ready
		.src_valid          (id_router_004_src_valid),                                            //          .valid
		.src_data           (id_router_004_src_data),                                             //          .data
		.src_channel        (id_router_004_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                       //          .endofpacket
	);

	nios2_system_id_router id_router_005 (
		.sink_ready         (switches_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (switches_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (switches_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (switches_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (switches_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                //       src.ready
		.src_valid          (id_router_005_src_valid),                                                //          .valid
		.src_data           (id_router_005_src_data),                                                 //          .data
		.src_channel        (id_router_005_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                           //          .endofpacket
	);

	nios2_system_id_router id_router_006 (
		.sink_ready         (key_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (key_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (key_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (key_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (key_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                           //       src.ready
		.src_valid          (id_router_006_src_valid),                                           //          .valid
		.src_data           (id_router_006_src_data),                                            //          .data
		.src_channel        (id_router_006_src_channel),                                         //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                   //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                      //          .endofpacket
	);

	nios2_system_id_router id_router_007 (
		.sink_ready         (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdcard_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                    //       src.ready
		.src_valid          (id_router_007_src_valid),                                                    //          .valid
		.src_data           (id_router_007_src_data),                                                     //          .data
		.src_channel        (id_router_007_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                               //          .endofpacket
	);

	nios2_system_id_router id_router_008 (
		.sink_ready         (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                                      // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                                                             //       src.ready
		.src_valid          (id_router_008_src_valid),                                                                                             //          .valid
		.src_data           (id_router_008_src_data),                                                                                              //          .data
		.src_channel        (id_router_008_src_channel),                                                                                           //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                                                                     //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                                                        //          .endofpacket
	);

	nios2_system_id_router id_router_009 (
		.sink_ready         (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ps2_0_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                           //       src.ready
		.src_valid          (id_router_009_src_valid),                                                           //          .valid
		.src_data           (id_router_009_src_data),                                                            //          .data
		.src_channel        (id_router_009_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                      //          .endofpacket
	);

	nios2_system_id_router id_router_010 (
		.sink_ready         (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (audio_0_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                               //       src.ready
		.src_valid          (id_router_010_src_valid),                                                               //          .valid
		.src_data           (id_router_010_src_data),                                                                //          .data
		.src_channel        (id_router_010_src_channel),                                                             //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                                          //          .endofpacket
	);

	nios2_system_id_router_011 id_router_011 (
		.sink_ready         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                                     //       src.ready
		.src_valid          (id_router_011_src_valid),                                                                     //          .valid
		.src_data           (id_router_011_src_data),                                                                      //          .data
		.src_channel        (id_router_011_src_channel),                                                                   //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                                             //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                                                //          .endofpacket
	);

	nios2_system_id_router_012 id_router_012 (
		.sink_ready         (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                           //       src.ready
		.src_valid          (id_router_012_src_valid),                                                           //          .valid
		.src_data           (id_router_012_src_data),                                                            //          .data
		.src_channel        (id_router_012_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                                      //          .endofpacket
	);

	nios2_system_id_router_012 id_router_013 (
		.sink_ready         (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (video_pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                         // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                                                //       src.ready
		.src_valid          (id_router_013_src_valid),                                                                                //          .valid
		.src_data           (id_router_013_src_data),                                                                                 //          .data
		.src_channel        (id_router_013_src_channel),                                                                              //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                                                        //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                                                           //          .endofpacket
	);

	nios2_system_id_router_012 id_router_014 (
		.sink_ready         (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (video_character_buffer_with_dma_0_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                                         // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                                                                                //       src.ready
		.src_valid          (id_router_014_src_valid),                                                                                                //          .valid
		.src_data           (id_router_014_src_data),                                                                                                 //          .data
		.src_channel        (id_router_014_src_channel),                                                                                              //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                                                                        //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                                                                           //          .endofpacket
	);

	nios2_system_id_router_011 id_router_015 (
		.sink_ready         (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (video_character_buffer_with_dma_0_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                                        // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                                                                               //       src.ready
		.src_valid          (id_router_015_src_valid),                                                                                               //          .valid
		.src_data           (id_router_015_src_data),                                                                                                //          .data
		.src_channel        (id_router_015_src_channel),                                                                                             //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                                                                       //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                                                                          //          .endofpacket
	);

	nios2_system_id_router_016 id_router_016 (
		.sink_ready         (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                                             //       src.ready
		.src_valid          (id_router_016_src_valid),                                                             //          .valid
		.src_data           (id_router_016_src_data),                                                              //          .data
		.src_channel        (id_router_016_src_channel),                                                           //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                                        //          .endofpacket
	);

	nios2_system_id_router_012 id_router_017 (
		.sink_ready         (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (audio_and_video_config_0_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                             // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                                                                    //       src.ready
		.src_valid          (id_router_017_src_valid),                                                                                    //          .valid
		.src_data           (id_router_017_src_data),                                                                                     //          .data
		.src_channel        (id_router_017_src_channel),                                                                                  //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                                                            //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                                                               //          .endofpacket
	);

	nios2_system_id_router_018 id_router_018 (
		.sink_ready         (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (usb_0_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                                                           //       src.ready
		.src_valid          (id_router_018_src_valid),                                                           //          .valid
		.src_data           (id_router_018_src_data),                                                            //          .data
		.src_channel        (id_router_018_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)                                                      //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (109),
		.ST_CHANNEL_W              (19),
		.VALID_WIDTH               (19),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clocks_sys_clk_clk),             //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (109),
		.ST_CHANNEL_W              (19),
		.VALID_WIDTH               (19),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (clocks_sys_clk_clk),                 //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_001_src_data),           //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (76),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.MAX_OUTSTANDING_RESPONSES (4),
		.PIPELINED                 (0),
		.ST_DATA_W                 (91),
		.ST_CHANNEL_W              (19),
		.VALID_WIDTH               (19),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16)
	) limiter_002 (
		.clk                    (clocks_sys_clk_clk),                 //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_002_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_002_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_002_src_data),           //          .data
		.cmd_sink_channel       (addr_router_002_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_002_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_002_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_002_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_002_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_002_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_002_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_002_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_002_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_002_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_002_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_002_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_002_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_002_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_002_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_002_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_002_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_002_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_002_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_002_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_002_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (69),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (91),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (57),
		.OUT_BURSTWRAP_H           (61),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (clocks_sys_clk_clk),                  //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_002_src_valid),          //     sink0.valid
		.sink0_data            (cmd_xbar_mux_002_src_data),           //          .data
		.sink0_channel         (cmd_xbar_mux_002_src_channel),        //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_002_src_startofpacket),  //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_002_src_endofpacket),    //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_002_src_ready),          //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (60),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.PKT_BURST_TYPE_H          (57),
		.PKT_BURST_TYPE_L          (56),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (82),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (47),
		.OUT_BURSTWRAP_H           (52),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_001 (
		.clk                   (clocks_sys_clk_clk),                      //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_002_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_002_src_data),              //          .data
		.sink0_channel         (width_adapter_002_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_002_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_002_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_002_src_ready),             //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (60),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.PKT_BURST_TYPE_H          (57),
		.PKT_BURST_TYPE_L          (56),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (82),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (47),
		.OUT_BURSTWRAP_H           (52),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_002 (
		.clk                   (clocks_sys_clk_clk),                      //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_003_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_003_src_data),              //          .data
		.sink0_channel         (width_adapter_003_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_003_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_003_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_003_src_ready),             //          .ready
		.source0_valid         (burst_adapter_002_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_002_source0_data),          //          .data
		.source0_channel       (burst_adapter_002_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_002_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_002_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_002_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (69),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (91),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (57),
		.OUT_BURSTWRAP_H           (61),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_003 (
		.clk                   (clocks_sys_clk_clk),                      //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_016_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_016_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_016_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_016_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_016_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_016_src_ready),              //          .ready
		.source0_valid         (burst_adapter_003_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_003_source0_data),          //          .data
		.source0_channel       (burst_adapter_003_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_003_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_003_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_003_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (1)
	) rst_controller (
		.reset_in0  (nios2_system_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1  (~reset_reset_n),                             // reset_in1.reset
		.clk        (clocks_sys_clk_clk),                         //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_req  (rst_controller_reset_out_reset_req),         //          .reset_req
		.reset_in2  (1'b0),                                       // (terminated)
		.reset_in3  (1'b0),                                       // (terminated)
		.reset_in4  (1'b0),                                       // (terminated)
		.reset_in5  (1'b0),                                       // (terminated)
		.reset_in6  (1'b0),                                       // (terminated)
		.reset_in7  (1'b0),                                       // (terminated)
		.reset_in8  (1'b0),                                       // (terminated)
		.reset_in9  (1'b0),                                       // (terminated)
		.reset_in10 (1'b0),                                       // (terminated)
		.reset_in11 (1'b0),                                       // (terminated)
		.reset_in12 (1'b0),                                       // (terminated)
		.reset_in13 (1'b0),                                       // (terminated)
		.reset_in14 (1'b0),                                       // (terminated)
		.reset_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_001 (
		.reset_in0  (nios2_system_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1  (~reset_reset_n),                             // reset_in1.reset
		.clk        (clk_clk),                                    //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),         // reset_out.reset
		.reset_req  (),                                           // (terminated)
		.reset_in2  (1'b0),                                       // (terminated)
		.reset_in3  (1'b0),                                       // (terminated)
		.reset_in4  (1'b0),                                       // (terminated)
		.reset_in5  (1'b0),                                       // (terminated)
		.reset_in6  (1'b0),                                       // (terminated)
		.reset_in7  (1'b0),                                       // (terminated)
		.reset_in8  (1'b0),                                       // (terminated)
		.reset_in9  (1'b0),                                       // (terminated)
		.reset_in10 (1'b0),                                       // (terminated)
		.reset_in11 (1'b0),                                       // (terminated)
		.reset_in12 (1'b0),                                       // (terminated)
		.reset_in13 (1'b0),                                       // (terminated)
		.reset_in14 (1'b0),                                       // (terminated)
		.reset_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_002 (
		.reset_in0  (nios2_system_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1  (~reset_reset_n),                             // reset_in1.reset
		.clk        (clocks_vga_clk_clk),                         //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset),         // reset_out.reset
		.reset_req  (),                                           // (terminated)
		.reset_in2  (1'b0),                                       // (terminated)
		.reset_in3  (1'b0),                                       // (terminated)
		.reset_in4  (1'b0),                                       // (terminated)
		.reset_in5  (1'b0),                                       // (terminated)
		.reset_in6  (1'b0),                                       // (terminated)
		.reset_in7  (1'b0),                                       // (terminated)
		.reset_in8  (1'b0),                                       // (terminated)
		.reset_in9  (1'b0),                                       // (terminated)
		.reset_in10 (1'b0),                                       // (terminated)
		.reset_in11 (1'b0),                                       // (terminated)
		.reset_in12 (1'b0),                                       // (terminated)
		.reset_in13 (1'b0),                                       // (terminated)
		.reset_in14 (1'b0),                                       // (terminated)
		.reset_in15 (1'b0)                                        // (terminated)
	);

	nios2_system_cmd_xbar_demux cmd_xbar_demux (
		.clk                 (clocks_sys_clk_clk),                 //        clk.clk
		.reset               (rst_controller_reset_out_reset),     //  clk_reset.reset
		.sink_ready          (limiter_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_cmd_src_channel),            //           .channel
		.sink_data           (limiter_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_src10_endofpacket)    //           .endofpacket
	);

	nios2_system_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (clocks_sys_clk_clk),                     //        clk.clk
		.reset               (rst_controller_reset_out_reset),         //  clk_reset.reset
		.sink_ready          (limiter_001_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_001_cmd_src_channel),            //           .channel
		.sink_data           (limiter_001_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_001_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_001_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_001_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //           .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //      src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //           .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //           .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //           .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //           .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //           .endofpacket
		.src12_ready         (cmd_xbar_demux_001_src12_ready),         //      src12.ready
		.src12_valid         (cmd_xbar_demux_001_src12_valid),         //           .valid
		.src12_data          (cmd_xbar_demux_001_src12_data),          //           .data
		.src12_channel       (cmd_xbar_demux_001_src12_channel),       //           .channel
		.src12_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //           .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_001_src12_endofpacket),   //           .endofpacket
		.src13_ready         (cmd_xbar_demux_001_src13_ready),         //      src13.ready
		.src13_valid         (cmd_xbar_demux_001_src13_valid),         //           .valid
		.src13_data          (cmd_xbar_demux_001_src13_data),          //           .data
		.src13_channel       (cmd_xbar_demux_001_src13_channel),       //           .channel
		.src13_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //           .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_001_src13_endofpacket),   //           .endofpacket
		.src14_ready         (cmd_xbar_demux_001_src14_ready),         //      src14.ready
		.src14_valid         (cmd_xbar_demux_001_src14_valid),         //           .valid
		.src14_data          (cmd_xbar_demux_001_src14_data),          //           .data
		.src14_channel       (cmd_xbar_demux_001_src14_channel),       //           .channel
		.src14_startofpacket (cmd_xbar_demux_001_src14_startofpacket), //           .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_001_src14_endofpacket),   //           .endofpacket
		.src15_ready         (cmd_xbar_demux_001_src15_ready),         //      src15.ready
		.src15_valid         (cmd_xbar_demux_001_src15_valid),         //           .valid
		.src15_data          (cmd_xbar_demux_001_src15_data),          //           .data
		.src15_channel       (cmd_xbar_demux_001_src15_channel),       //           .channel
		.src15_startofpacket (cmd_xbar_demux_001_src15_startofpacket), //           .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_001_src15_endofpacket),   //           .endofpacket
		.src16_ready         (cmd_xbar_demux_001_src16_ready),         //      src16.ready
		.src16_valid         (cmd_xbar_demux_001_src16_valid),         //           .valid
		.src16_data          (cmd_xbar_demux_001_src16_data),          //           .data
		.src16_channel       (cmd_xbar_demux_001_src16_channel),       //           .channel
		.src16_startofpacket (cmd_xbar_demux_001_src16_startofpacket), //           .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_001_src16_endofpacket),   //           .endofpacket
		.src17_ready         (cmd_xbar_demux_001_src17_ready),         //      src17.ready
		.src17_valid         (cmd_xbar_demux_001_src17_valid),         //           .valid
		.src17_data          (cmd_xbar_demux_001_src17_data),          //           .data
		.src17_channel       (cmd_xbar_demux_001_src17_channel),       //           .channel
		.src17_startofpacket (cmd_xbar_demux_001_src17_startofpacket), //           .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_001_src17_endofpacket),   //           .endofpacket
		.src18_ready         (cmd_xbar_demux_001_src18_ready),         //      src18.ready
		.src18_valid         (cmd_xbar_demux_001_src18_valid),         //           .valid
		.src18_data          (cmd_xbar_demux_001_src18_data),          //           .data
		.src18_channel       (cmd_xbar_demux_001_src18_channel),       //           .channel
		.src18_startofpacket (cmd_xbar_demux_001_src18_startofpacket), //           .startofpacket
		.src18_endofpacket   (cmd_xbar_demux_001_src18_endofpacket)    //           .endofpacket
	);

	nios2_system_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (clocks_sys_clk_clk),                    //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_002_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_002_cmd_src_channel),           //           .channel
		.sink_data          (limiter_002_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_002_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_002_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_002_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_002_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_002_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_002_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_002_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_002_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_002_src1_endofpacket)    //           .endofpacket
	);

	nios2_system_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios2_system_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	nios2_system_cmd_xbar_mux_002 cmd_xbar_mux_002 (
		.clk                 (clocks_sys_clk_clk),                  //       clk.clk
		.reset               (rst_controller_reset_out_reset),      // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),          //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),          //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),           //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),        //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),  //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),    //          .endofpacket
		.sink0_ready         (width_adapter_src_ready),             //     sink0.ready
		.sink0_valid         (width_adapter_src_valid),             //          .valid
		.sink0_channel       (width_adapter_src_channel),           //          .channel
		.sink0_data          (width_adapter_src_data),              //          .data
		.sink0_startofpacket (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (width_adapter_src_endofpacket),       //          .endofpacket
		.sink1_ready         (width_adapter_001_src_ready),         //     sink1.ready
		.sink1_valid         (width_adapter_001_src_valid),         //          .valid
		.sink1_channel       (width_adapter_001_src_channel),       //          .channel
		.sink1_data          (width_adapter_001_src_data),          //          .data
		.sink1_startofpacket (width_adapter_001_src_startofpacket), //          .startofpacket
		.sink1_endofpacket   (width_adapter_001_src_endofpacket)    //          .endofpacket
	);

	nios2_system_cmd_xbar_mux cmd_xbar_mux_003 (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src3_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src3_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src3_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src3_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src3_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src3_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src3_endofpacket)    //          .endofpacket
	);

	nios2_system_cmd_xbar_mux cmd_xbar_mux_004 (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_004_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_004_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_004_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_004_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_004_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_004_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src4_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src4_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src4_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src4_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src4_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src4_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src4_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src4_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src4_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src4_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src4_endofpacket)    //          .endofpacket
	);

	nios2_system_cmd_xbar_mux cmd_xbar_mux_005 (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_005_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_005_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_005_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_005_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_005_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_005_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src5_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src5_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src5_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src5_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src5_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src5_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src5_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src5_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src5_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src5_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src5_endofpacket)    //          .endofpacket
	);

	nios2_system_cmd_xbar_mux cmd_xbar_mux_006 (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_006_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_006_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_006_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_006_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_006_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_006_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src6_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src6_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src6_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src6_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src6_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src6_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src6_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src6_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src6_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src6_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src6_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src6_endofpacket)    //          .endofpacket
	);

	nios2_system_cmd_xbar_mux cmd_xbar_mux_007 (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_007_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_007_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_007_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_007_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_007_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_007_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src7_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src7_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src7_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src7_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src7_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src7_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src7_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src7_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src7_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src7_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src7_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src7_endofpacket)    //          .endofpacket
	);

	nios2_system_cmd_xbar_mux cmd_xbar_mux_008 (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_008_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_008_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_008_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_008_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_008_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_008_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src8_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src8_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src8_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src8_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src8_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src8_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src8_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src8_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src8_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src8_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src8_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src8_endofpacket)    //          .endofpacket
	);

	nios2_system_cmd_xbar_mux cmd_xbar_mux_009 (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_009_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_009_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_009_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_009_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_009_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_009_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src9_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src9_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src9_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src9_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src9_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src9_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src9_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src9_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src9_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src9_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src9_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src9_endofpacket)    //          .endofpacket
	);

	nios2_system_cmd_xbar_mux cmd_xbar_mux_010 (
		.clk                 (clocks_sys_clk_clk),                     //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.src_ready           (cmd_xbar_mux_010_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_010_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_010_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_010_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_010_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_010_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src10_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src10_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src10_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src10_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src10_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src10_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src10_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src10_endofpacket)    //          .endofpacket
	);

	nios2_system_cmd_xbar_mux_002 cmd_xbar_mux_016 (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_016_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_016_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_016_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_016_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_016_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_016_src_endofpacket),      //          .endofpacket
		.sink0_ready         (width_adapter_004_src_ready),           //     sink0.ready
		.sink0_valid         (width_adapter_004_src_valid),           //          .valid
		.sink0_channel       (width_adapter_004_src_channel),         //          .channel
		.sink0_data          (width_adapter_004_src_data),            //          .data
		.sink0_startofpacket (width_adapter_004_src_startofpacket),   //          .startofpacket
		.sink0_endofpacket   (width_adapter_004_src_endofpacket),     //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios2_system_cmd_xbar_mux cmd_xbar_mux_018 (
		.clk                 (clocks_sys_clk_clk),                     //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.src_ready           (cmd_xbar_mux_018_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_018_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_018_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_018_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_018_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_018_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src18_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src18_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src18_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src18_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src18_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src18_endofpacket),   //          .endofpacket
		.sink1_ready         (width_adapter_005_src_ready),            //     sink1.ready
		.sink1_valid         (width_adapter_005_src_valid),            //          .valid
		.sink1_channel       (width_adapter_005_src_channel),          //          .channel
		.sink1_data          (width_adapter_005_src_data),             //          .data
		.sink1_startofpacket (width_adapter_005_src_startofpacket),    //          .startofpacket
		.sink1_endofpacket   (width_adapter_005_src_endofpacket)       //          .endofpacket
	);

	nios2_system_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clocks_sys_clk_clk),                //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	nios2_system_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	nios2_system_rsp_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	nios2_system_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	nios2_system_rsp_xbar_demux rsp_xbar_demux_004 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_004_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_004_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_004_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_004_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_004_src1_endofpacket)    //          .endofpacket
	);

	nios2_system_rsp_xbar_demux rsp_xbar_demux_005 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_005_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_005_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_005_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_005_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_005_src1_endofpacket)    //          .endofpacket
	);

	nios2_system_rsp_xbar_demux rsp_xbar_demux_006 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_006_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_006_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_006_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_006_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_006_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_006_src1_endofpacket)    //          .endofpacket
	);

	nios2_system_rsp_xbar_demux rsp_xbar_demux_007 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_007_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_007_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_007_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_007_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_007_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_007_src1_endofpacket)    //          .endofpacket
	);

	nios2_system_rsp_xbar_demux rsp_xbar_demux_008 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_008_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_008_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_008_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_008_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_008_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_008_src1_endofpacket)    //          .endofpacket
	);

	nios2_system_rsp_xbar_demux rsp_xbar_demux_009 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_009_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_009_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_009_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_009_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_009_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_009_src1_endofpacket)    //          .endofpacket
	);

	nios2_system_rsp_xbar_demux rsp_xbar_demux_010 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_010_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_010_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_010_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_010_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_010_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_010_src1_endofpacket)    //          .endofpacket
	);

	nios2_system_rsp_xbar_demux_011 rsp_xbar_demux_011 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	nios2_system_rsp_xbar_demux_012 rsp_xbar_demux_012 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	nios2_system_rsp_xbar_demux_012 rsp_xbar_demux_013 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	nios2_system_rsp_xbar_demux_012 rsp_xbar_demux_014 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	nios2_system_rsp_xbar_demux_011 rsp_xbar_demux_015 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	nios2_system_rsp_xbar_demux_002 rsp_xbar_demux_016 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_016_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_016_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_016_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_016_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_016_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_016_src1_endofpacket)    //          .endofpacket
	);

	nios2_system_rsp_xbar_demux_012 rsp_xbar_demux_017 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	nios2_system_rsp_xbar_demux rsp_xbar_demux_018 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_018_src_ready),               //      sink.ready
		.sink_channel       (id_router_018_src_channel),             //          .channel
		.sink_data          (id_router_018_src_data),                //          .data
		.sink_startofpacket (id_router_018_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_018_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_018_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_018_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_018_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_018_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_018_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_018_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_018_src1_endofpacket)    //          .endofpacket
	);

	nios2_system_rsp_xbar_mux rsp_xbar_mux (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid            (rsp_xbar_mux_src_valid),                //          .valid
		.src_data             (rsp_xbar_mux_src_data),                 //          .data
		.src_channel          (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket    (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready          (width_adapter_006_src_ready),           //     sink2.ready
		.sink2_valid          (width_adapter_006_src_valid),           //          .valid
		.sink2_channel        (width_adapter_006_src_channel),         //          .channel
		.sink2_data           (width_adapter_006_src_data),            //          .data
		.sink2_startofpacket  (width_adapter_006_src_startofpacket),   //          .startofpacket
		.sink2_endofpacket    (width_adapter_006_src_endofpacket),     //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	nios2_system_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (width_adapter_007_src_ready),           //     sink2.ready
		.sink2_valid          (width_adapter_007_src_valid),           //          .valid
		.sink2_channel        (width_adapter_007_src_channel),         //          .channel
		.sink2_data           (width_adapter_007_src_data),            //          .data
		.sink2_startofpacket  (width_adapter_007_src_startofpacket),   //          .startofpacket
		.sink2_endofpacket    (width_adapter_007_src_endofpacket),     //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src1_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src1_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src1_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src1_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src1_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src1_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src1_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src1_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src1_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src1_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src1_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src1_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src1_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src1_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src1_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src1_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src1_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src1_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src1_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src1_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src1_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src1_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src1_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src1_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src1_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src1_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src1_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src1_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src1_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src1_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src1_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src1_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src1_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src1_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src1_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src1_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src1_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src1_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src1_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src1_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src1_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src1_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src1_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src1_endofpacket),   //          .endofpacket
		.sink11_ready         (width_adapter_008_src_ready),           //    sink11.ready
		.sink11_valid         (width_adapter_008_src_valid),           //          .valid
		.sink11_channel       (width_adapter_008_src_channel),         //          .channel
		.sink11_data          (width_adapter_008_src_data),            //          .data
		.sink11_startofpacket (width_adapter_008_src_startofpacket),   //          .startofpacket
		.sink11_endofpacket   (width_adapter_008_src_endofpacket),     //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_014_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (width_adapter_009_src_ready),           //    sink15.ready
		.sink15_valid         (width_adapter_009_src_valid),           //          .valid
		.sink15_channel       (width_adapter_009_src_channel),         //          .channel
		.sink15_data          (width_adapter_009_src_data),            //          .data
		.sink15_startofpacket (width_adapter_009_src_startofpacket),   //          .startofpacket
		.sink15_endofpacket   (width_adapter_009_src_endofpacket),     //          .endofpacket
		.sink16_ready         (width_adapter_010_src_ready),           //    sink16.ready
		.sink16_valid         (width_adapter_010_src_valid),           //          .valid
		.sink16_channel       (width_adapter_010_src_channel),         //          .channel
		.sink16_data          (width_adapter_010_src_data),            //          .data
		.sink16_startofpacket (width_adapter_010_src_startofpacket),   //          .startofpacket
		.sink16_endofpacket   (width_adapter_010_src_endofpacket),     //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_017_src0_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_017_src0_endofpacket),   //          .endofpacket
		.sink18_ready         (rsp_xbar_demux_018_src0_ready),         //    sink18.ready
		.sink18_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.sink18_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.sink18_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.sink18_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.sink18_endofpacket   (rsp_xbar_demux_018_src0_endofpacket)    //          .endofpacket
	);

	nios2_system_rsp_xbar_mux_002 rsp_xbar_mux_002 (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_002_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_002_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_016_src1_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_016_src1_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_016_src1_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_016_src1_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_016_src1_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_016_src1_endofpacket),   //          .endofpacket
		.sink1_ready         (width_adapter_011_src_ready),           //     sink1.ready
		.sink1_valid         (width_adapter_011_src_valid),           //          .valid
		.sink1_channel       (width_adapter_011_src_channel),         //          .channel
		.sink1_data          (width_adapter_011_src_data),            //          .data
		.sink1_startofpacket (width_adapter_011_src_startofpacket),   //          .startofpacket
		.sink1_endofpacket   (width_adapter_011_src_endofpacket)      //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (108),
		.IN_PKT_RESPONSE_STATUS_L      (107),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (109),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (90),
		.OUT_PKT_RESPONSE_STATUS_L     (89),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (91),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter (
		.clk                  (clocks_sys_clk_clk),                //       clk.clk
		.reset                (rst_controller_reset_out_reset),    // clk_reset.reset
		.in_valid             (cmd_xbar_demux_src2_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_src2_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_src2_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_src2_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_src2_ready),         //          .ready
		.in_data              (cmd_xbar_demux_src2_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_src_data),            //          .data
		.out_channel          (width_adapter_src_channel),         //          .channel
		.out_valid            (width_adapter_src_valid),           //          .valid
		.out_ready            (width_adapter_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                             // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (108),
		.IN_PKT_RESPONSE_STATUS_L      (107),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (109),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (90),
		.OUT_PKT_RESPONSE_STATUS_L     (89),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (91),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_001 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src2_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src2_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src2_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src2_data),          //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_001_src_data),            //          .data
		.out_channel          (width_adapter_001_src_channel),         //          .channel
		.out_valid            (width_adapter_001_src_valid),           //          .valid
		.out_ready            (width_adapter_001_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (108),
		.IN_PKT_RESPONSE_STATUS_L      (107),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (109),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (49),
		.OUT_PKT_BYTE_CNT_L            (47),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_PKT_BURST_SIZE_H          (55),
		.OUT_PKT_BURST_SIZE_L          (53),
		.OUT_PKT_RESPONSE_STATUS_H     (81),
		.OUT_PKT_RESPONSE_STATUS_L     (80),
		.OUT_PKT_TRANS_EXCLUSIVE       (46),
		.OUT_PKT_BURST_TYPE_H          (57),
		.OUT_PKT_BURST_TYPE_L          (56),
		.OUT_ST_DATA_W                 (82),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_002 (
		.clk                  (clocks_sys_clk_clk),                     //       clk.clk
		.reset                (rst_controller_reset_out_reset),         // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src11_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src11_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src11_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src11_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src11_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src11_data),          //          .data
		.out_endofpacket      (width_adapter_002_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_002_src_data),             //          .data
		.out_channel          (width_adapter_002_src_channel),          //          .channel
		.out_valid            (width_adapter_002_src_valid),            //          .valid
		.out_ready            (width_adapter_002_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_002_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                                  // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (108),
		.IN_PKT_RESPONSE_STATUS_L      (107),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (109),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (49),
		.OUT_PKT_BYTE_CNT_L            (47),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_PKT_BURST_SIZE_H          (55),
		.OUT_PKT_BURST_SIZE_L          (53),
		.OUT_PKT_RESPONSE_STATUS_H     (81),
		.OUT_PKT_RESPONSE_STATUS_L     (80),
		.OUT_PKT_TRANS_EXCLUSIVE       (46),
		.OUT_PKT_BURST_TYPE_H          (57),
		.OUT_PKT_BURST_TYPE_L          (56),
		.OUT_ST_DATA_W                 (82),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_003 (
		.clk                  (clocks_sys_clk_clk),                     //       clk.clk
		.reset                (rst_controller_reset_out_reset),         // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src15_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src15_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src15_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src15_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src15_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src15_data),          //          .data
		.out_endofpacket      (width_adapter_003_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_003_src_data),             //          .data
		.out_channel          (width_adapter_003_src_channel),          //          .channel
		.out_valid            (width_adapter_003_src_valid),            //          .valid
		.out_ready            (width_adapter_003_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_003_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                                  // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (108),
		.IN_PKT_RESPONSE_STATUS_L      (107),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (109),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (90),
		.OUT_PKT_RESPONSE_STATUS_L     (89),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (91),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_004 (
		.clk                  (clocks_sys_clk_clk),                     //       clk.clk
		.reset                (rst_controller_reset_out_reset),         // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src16_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src16_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src16_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src16_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src16_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src16_data),          //          .data
		.out_endofpacket      (width_adapter_004_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_004_src_data),             //          .data
		.out_channel          (width_adapter_004_src_channel),          //          .channel
		.out_valid            (width_adapter_004_src_valid),            //          .valid
		.out_ready            (width_adapter_004_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_004_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                                  // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (90),
		.IN_PKT_RESPONSE_STATUS_L      (89),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (91),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (108),
		.OUT_PKT_RESPONSE_STATUS_L     (107),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (109),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_005 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_002_src1_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_002_src1_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_002_src1_ready),         //          .ready
		.in_data              (cmd_xbar_demux_002_src1_data),          //          .data
		.out_endofpacket      (width_adapter_005_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_005_src_data),            //          .data
		.out_channel          (width_adapter_005_src_channel),         //          .channel
		.out_valid            (width_adapter_005_src_valid),           //          .valid
		.out_ready            (width_adapter_005_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_005_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (90),
		.IN_PKT_RESPONSE_STATUS_L      (89),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (91),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (108),
		.OUT_PKT_RESPONSE_STATUS_L     (107),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (109),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_006 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_002_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_002_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_002_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_002_src0_data),          //          .data
		.out_endofpacket      (width_adapter_006_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_006_src_data),            //          .data
		.out_channel          (width_adapter_006_src_channel),         //          .channel
		.out_valid            (width_adapter_006_src_valid),           //          .valid
		.out_ready            (width_adapter_006_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_006_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (90),
		.IN_PKT_RESPONSE_STATUS_L      (89),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (91),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (108),
		.OUT_PKT_RESPONSE_STATUS_L     (107),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (109),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_007 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_002_src1_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_002_src1_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_002_src1_ready),         //          .ready
		.in_data              (rsp_xbar_demux_002_src1_data),          //          .data
		.out_endofpacket      (width_adapter_007_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_007_src_data),            //          .data
		.out_channel          (width_adapter_007_src_channel),         //          .channel
		.out_valid            (width_adapter_007_src_valid),           //          .valid
		.out_ready            (width_adapter_007_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_007_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (49),
		.IN_PKT_BYTE_CNT_L             (47),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (52),
		.IN_PKT_BURSTWRAP_L            (50),
		.IN_PKT_BURST_SIZE_H           (55),
		.IN_PKT_BURST_SIZE_L           (53),
		.IN_PKT_RESPONSE_STATUS_H      (81),
		.IN_PKT_RESPONSE_STATUS_L      (80),
		.IN_PKT_TRANS_EXCLUSIVE        (46),
		.IN_PKT_BURST_TYPE_H           (57),
		.IN_PKT_BURST_TYPE_L           (56),
		.IN_ST_DATA_W                  (82),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (108),
		.OUT_PKT_RESPONSE_STATUS_L     (107),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (109),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_008 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_011_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_011_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_011_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_011_src0_data),          //          .data
		.out_endofpacket      (width_adapter_008_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_008_src_data),            //          .data
		.out_channel          (width_adapter_008_src_channel),         //          .channel
		.out_valid            (width_adapter_008_src_valid),           //          .valid
		.out_ready            (width_adapter_008_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_008_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (49),
		.IN_PKT_BYTE_CNT_L             (47),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (52),
		.IN_PKT_BURSTWRAP_L            (50),
		.IN_PKT_BURST_SIZE_H           (55),
		.IN_PKT_BURST_SIZE_L           (53),
		.IN_PKT_RESPONSE_STATUS_H      (81),
		.IN_PKT_RESPONSE_STATUS_L      (80),
		.IN_PKT_TRANS_EXCLUSIVE        (46),
		.IN_PKT_BURST_TYPE_H           (57),
		.IN_PKT_BURST_TYPE_L           (56),
		.IN_ST_DATA_W                  (82),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (108),
		.OUT_PKT_RESPONSE_STATUS_L     (107),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (109),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_009 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_015_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_015_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_015_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_015_src0_data),          //          .data
		.out_endofpacket      (width_adapter_009_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_009_src_data),            //          .data
		.out_channel          (width_adapter_009_src_channel),         //          .channel
		.out_valid            (width_adapter_009_src_valid),           //          .valid
		.out_ready            (width_adapter_009_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_009_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (90),
		.IN_PKT_RESPONSE_STATUS_L      (89),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (91),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (108),
		.OUT_PKT_RESPONSE_STATUS_L     (107),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (109),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_010 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_016_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_016_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_016_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_016_src0_data),          //          .data
		.out_endofpacket      (width_adapter_010_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_010_src_data),            //          .data
		.out_channel          (width_adapter_010_src_channel),         //          .channel
		.out_valid            (width_adapter_010_src_valid),           //          .valid
		.out_ready            (width_adapter_010_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_010_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (108),
		.IN_PKT_RESPONSE_STATUS_L      (107),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (109),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (90),
		.OUT_PKT_RESPONSE_STATUS_L     (89),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (91),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_011 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_018_src1_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_018_src1_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_018_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_018_src1_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_018_src1_ready),         //          .ready
		.in_data              (rsp_xbar_demux_018_src1_data),          //          .data
		.out_endofpacket      (width_adapter_011_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_011_src_data),            //          .data
		.out_channel          (width_adapter_011_src_channel),         //          .channel
		.out_valid            (width_adapter_011_src_valid),           //          .valid
		.out_ready            (width_adapter_011_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_011_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	nios2_system_irq_mapper irq_mapper (
		.clk           (clocks_sys_clk_clk),             //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (nios2_system_d_irq_irq)          //    sender.irq
	);

endmodule
